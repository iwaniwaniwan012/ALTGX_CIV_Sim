-- megafunction wizard: %ALTGX_RECONFIG%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: alt_c3gxb_reconfig 

-- ============================================================
-- File Name: ALTGX_RECONFIG_CIV.vhd
-- Megafunction Name(s):
-- 			alt_c3gxb_reconfig
--
-- Simulation Library Files(s):
-- 			altera_mf;lpm
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 21.1.0 Build 842 10/21/2021 SJ Lite Edition
-- ************************************************************


--Copyright (C) 2021  Intel Corporation. All rights reserved.
--Your use of Intel Corporation's design tools, logic functions 
--and other software and tools, and any partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Intel Program License 
--Subscription Agreement, the Intel Quartus Prime License Agreement,
--the Intel FPGA IP License Agreement, or other applicable license
--agreement, including, without limitation, that your use is for
--the sole purpose of programming logic devices manufactured by
--Intel and sold by Intel or its authorized distributors.  Please
--refer to the applicable agreement for further details, at
--https://fpgasoftware.intel.com/eula.


--alt_c3gxb_reconfig CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone IV GX" ENABLE_BUF_CAL="TRUE" ENABLE_ILLEGAL_MODE_CHECK="TRUE" ENABLE_SELF_RECOVERY="TRUE" MIF_ADDRESS_WIDTH=6 NUMBER_OF_CHANNELS=1 NUMBER_OF_RECONFIG_PORTS=1 RECONFIG_FROMGXB_WIDTH=5 RECONFIG_TOGXB_WIDTH=4 busy channel_reconfig_done error reconfig_address_en reconfig_address_out reconfig_clk reconfig_data reconfig_fromgxb reconfig_mode_sel reconfig_reset reconfig_togxb write_all
--VERSION_BEGIN 21.1 cbx_alt_c3gxb_reconfig 2021:10:21:11:02:24:SJ cbx_alt_cal 2021:10:21:11:02:24:SJ cbx_alt_dprio 2021:10:21:11:02:24:SJ cbx_altera_syncram_nd_impl 2021:10:21:11:02:24:SJ cbx_altsyncram 2021:10:21:11:02:24:SJ cbx_cycloneii 2021:10:21:11:02:24:SJ cbx_lpm_add_sub 2021:10:21:11:02:24:SJ cbx_lpm_compare 2021:10:21:11:02:24:SJ cbx_lpm_counter 2021:10:21:11:02:24:SJ cbx_lpm_decode 2021:10:21:11:02:24:SJ cbx_lpm_mux 2021:10:21:11:02:24:SJ cbx_lpm_shiftreg 2021:10:21:11:02:24:SJ cbx_mgl 2021:10:21:11:11:47:SJ cbx_nadder 2021:10:21:11:02:24:SJ cbx_stratix 2021:10:21:11:02:24:SJ cbx_stratixii 2021:10:21:11:02:24:SJ cbx_stratixiii 2021:10:21:11:02:24:SJ cbx_stratixv 2021:10:21:11:02:24:SJ cbx_util_mgl 2021:10:21:11:02:24:SJ  VERSION_END


--alt_dprio address_width=16 CBX_AUTO_BLACKBOX="ALL" device_family="Cyclone IV GX" quad_address_width=9 address busy datain dataout dpclk dpriodisable dprioin dprioload dprioout quad_address rden reset status_out wren wren_data
--VERSION_BEGIN 21.1 cbx_alt_dprio 2021:10:21:11:02:24:SJ cbx_cycloneii 2021:10:21:11:02:24:SJ cbx_lpm_add_sub 2021:10:21:11:02:24:SJ cbx_lpm_compare 2021:10:21:11:02:24:SJ cbx_lpm_counter 2021:10:21:11:02:24:SJ cbx_lpm_decode 2021:10:21:11:02:24:SJ cbx_lpm_shiftreg 2021:10:21:11:02:24:SJ cbx_mgl 2021:10:21:11:11:47:SJ cbx_nadder 2021:10:21:11:02:24:SJ cbx_stratix 2021:10:21:11:02:24:SJ cbx_stratixii 2021:10:21:11:02:24:SJ  VERSION_END

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = lpm_compare 3 lpm_counter 1 lpm_decode 1 lut 1 reg 102 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  ALTGX_RECONFIG_CIV_alt_dprio_q9l IS 
	 PORT 
	 ( 
		 address	:	IN  STD_LOGIC_VECTOR (15 DOWNTO 0);
		 busy	:	OUT  STD_LOGIC;
		 datain	:	IN  STD_LOGIC_VECTOR (15 DOWNTO 0) := (OTHERS => '0');
		 dataout	:	OUT  STD_LOGIC_VECTOR (15 DOWNTO 0);
		 dpclk	:	IN  STD_LOGIC;
		 dpriodisable	:	OUT  STD_LOGIC;
		 dprioin	:	OUT  STD_LOGIC;
		 dprioload	:	OUT  STD_LOGIC;
		 dprioout	:	IN  STD_LOGIC;
		 quad_address	:	IN  STD_LOGIC_VECTOR (8 DOWNTO 0);
		 rden	:	IN  STD_LOGIC := '0';
		 reset	:	IN  STD_LOGIC := '0';
		 status_out	:	OUT  STD_LOGIC_VECTOR (3 DOWNTO 0);
		 wren	:	IN  STD_LOGIC := '0';
		 wren_data	:	IN  STD_LOGIC := '0'
	 ); 
 END ALTGX_RECONFIG_CIV_alt_dprio_q9l;

 ARCHITECTURE RTL OF ALTGX_RECONFIG_CIV_alt_dprio_q9l IS

	 ATTRIBUTE synthesis_clearbox : natural;
	 ATTRIBUTE synthesis_clearbox OF RTL : ARCHITECTURE IS 2;
	 ATTRIBUTE ALTERA_ATTRIBUTE : string;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF RTL : ARCHITECTURE IS "{-to addr_shift_reg[31]} DPRIO_INTERFACE_REG=ON;{-to wr_out_data_shift_reg[31]} DPRIO_INTERFACE_REG=ON;{-to rd_out_data_shift_reg[13]} DPRIO_INTERFACE_REG=ON;{-to in_data_shift_reg[0]} DPRIO_INTERFACE_REG=ON;{-to startup_cntr[0]} DPRIO_INTERFACE_REG=ON;{-to startup_cntr[1]} DPRIO_INTERFACE_REG=ON;{-to startup_cntr[2]} DPRIO_INTERFACE_REG=ON";

	 SIGNAL	 wire_addr_shift_reg_d	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL	 wire_addr_shift_reg_asdata	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL	 addr_shift_reg	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF addr_shift_reg : SIGNAL IS "PRESERVE_REGISTER=ON;POWER_UP_LEVEL=LOW";

	 SIGNAL  wire_addr_shift_reg_w_q_range862w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 in_data_shift_reg	:	STD_LOGIC_VECTOR(15 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF in_data_shift_reg : SIGNAL IS "PRESERVE_REGISTER=ON;POWER_UP_LEVEL=LOW";

	 SIGNAL	 wire_rd_out_data_shift_reg_d	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL	 wire_rd_out_data_shift_reg_asdata	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL	 rd_out_data_shift_reg	:	STD_LOGIC_VECTOR(15 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF rd_out_data_shift_reg : SIGNAL IS "PRESERVE_REGISTER=ON;POWER_UP_LEVEL=LOW";

	 SIGNAL  wire_rd_out_data_shift_reg_w_q_range1038w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 wire_startup_cntr_d	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL	 startup_cntr	:	STD_LOGIC_VECTOR(2 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF startup_cntr : SIGNAL IS "PRESERVE_REGISTER=ON;POWER_UP_LEVEL=LOW";

	 SIGNAL	 wire_startup_cntr_ena	:	STD_LOGIC_VECTOR(2 DOWNTO 0);
	 SIGNAL  wire_startup_cntr_w_lg_w_q_range1103w1106w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_startup_cntr_w_lg_w_q_range1107w1113w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_startup_cntr_w_lg_w_q_range1107w1116w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_startup_cntr_w_lg_w_q_range1099w1100w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_startup_cntr_w_lg_w_q_range1099w1115w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_startup_cntr_w_lg_w_q_range1099w1104w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_startup_cntr_w_lg_w_q_range1107w1108w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_startup_cntr_w_q_range1099w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_startup_cntr_w_q_range1103w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_startup_cntr_w_q_range1107w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 state_mc_reg	:	STD_LOGIC_VECTOR(2 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF state_mc_reg : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL  wire_state_mc_reg_w_q_range692w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_state_mc_reg_w_q_range711w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_state_mc_reg_w_q_range727w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 wire_wr_out_data_shift_reg_d	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL	 wire_wr_out_data_shift_reg_asdata	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL	 wr_out_data_shift_reg	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF wr_out_data_shift_reg : SIGNAL IS "PRESERVE_REGISTER=ON;POWER_UP_LEVEL=LOW";

	 SIGNAL  wire_wr_out_data_shift_reg_w_q_range973w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_pre_amble_cmpr_w_lg_w_lg_agb860w1037w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_pre_amble_cmpr_w_lg_w_lg_agb860w972w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_pre_amble_cmpr_w_lg_agb860w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_pre_amble_cmpr_aeb	:	STD_LOGIC;
	 SIGNAL  wire_pre_amble_cmpr_agb	:	STD_LOGIC;
	 SIGNAL  wire_pre_amble_cmpr_datab	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_rd_data_output_cmpr_ageb	:	STD_LOGIC;
	 SIGNAL  wire_rd_data_output_cmpr_alb	:	STD_LOGIC;
	 SIGNAL  wire_rd_data_output_cmpr_datab	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_state_mc_cmpr_aeb	:	STD_LOGIC;
	 SIGNAL  wire_state_mc_cmpr_datab	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_state_mc_counter_cnt_en	:	STD_LOGIC;
	 SIGNAL  wire_dprio_w_lg_write_state677w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_state_mc_counter_q	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_state_mc_decode_eq	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL	wire_dprioin_mux_dataout	:	STD_LOGIC;
	 SIGNAL  wire_dprio_w_lg_w_lg_w_lg_s0_to_0694w695w696w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_w_lg_s1_to_0713w714w715w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_w_lg_s2_to_0729w730w731w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_w_lg_wren683w706w719w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_w_lg_wren683w706w707w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_w_lg_wr_addr_state859w863w864w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_rd_data_output_state1039w1040w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_wr_data_state974w975w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_s0_to_0694w695w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_s1_to_0713w714w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_s2_to_0729w730w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_wren683w706w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_wren683w684w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_wren683w701w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_w_lg_w_lg_rden1095w1096w1097w1098w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_wr_addr_state859w863w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_idle_state720w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_idle_state702w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_idle_state709w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_idle_state686w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_idle_state723w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_rd_data_output_state1039w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_wr_data_state974w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_s0_to_0694w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_s0_to_1693w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_s1_to_0713w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_s1_to_1712w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_s2_to_0729w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_s2_to_1728w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_startup_done1093w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_startup_idle1094w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_wren683w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_wren_data705w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_w_lg_rden1095w1096w1097w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_rden681w682w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_rden1095w1096w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_rden681w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_rden1095w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_rdinc718w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_rdinc700w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_s0_to_1697w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_s1_to_1716w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_s2_to_1732w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_wr_addr_state859w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_wren708w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_wren685w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_wren722w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  busy_state :	STD_LOGIC;
	 SIGNAL  idle_state :	STD_LOGIC;
	 SIGNAL  rd_addr_done :	STD_LOGIC;
	 SIGNAL  rd_addr_state :	STD_LOGIC;
	 SIGNAL  rd_data_done :	STD_LOGIC;
	 SIGNAL  rd_data_input_state :	STD_LOGIC;
	 SIGNAL  rd_data_output_state :	STD_LOGIC;
	 SIGNAL  rd_data_state :	STD_LOGIC;
	 SIGNAL  rdinc	:	STD_LOGIC;
	 SIGNAL  read_state :	STD_LOGIC;
	 SIGNAL  s0_to_0 :	STD_LOGIC;
	 SIGNAL  s0_to_1 :	STD_LOGIC;
	 SIGNAL  s1_to_0 :	STD_LOGIC;
	 SIGNAL  s1_to_1 :	STD_LOGIC;
	 SIGNAL  s2_to_0 :	STD_LOGIC;
	 SIGNAL  s2_to_1 :	STD_LOGIC;
	 SIGNAL  startup_done :	STD_LOGIC;
	 SIGNAL  startup_idle :	STD_LOGIC;
	 SIGNAL  wr_addr_done :	STD_LOGIC;
	 SIGNAL  wr_addr_state :	STD_LOGIC;
	 SIGNAL  wr_data_done :	STD_LOGIC;
	 SIGNAL  wr_data_state :	STD_LOGIC;
	 SIGNAL  write_state :	STD_LOGIC;
	 COMPONENT  lpm_compare
	 GENERIC 
	 (
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "UNSIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_compare"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		aeb	:	OUT STD_LOGIC;
		agb	:	OUT STD_LOGIC;
		ageb	:	OUT STD_LOGIC;
		alb	:	OUT STD_LOGIC;
		aleb	:	OUT STD_LOGIC;
		aneb	:	OUT STD_LOGIC;
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_counter
	 GENERIC 
	 (
		lpm_avalue	:	STRING := "0";
		lpm_direction	:	STRING := "DEFAULT";
		lpm_modulus	:	NATURAL := 0;
		lpm_port_updown	:	STRING := "PORT_CONNECTIVITY";
		lpm_pvalue	:	STRING := "0";
		lpm_svalue	:	STRING := "0";
		lpm_width	:	NATURAL;
		lpm_type	:	STRING := "lpm_counter"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		aload	:	IN STD_LOGIC := '0';
		aset	:	IN STD_LOGIC := '0';
		cin	:	IN STD_LOGIC := '1';
		clk_en	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC;
		cnt_en	:	IN STD_LOGIC := '1';
		cout	:	OUT STD_LOGIC;
		data	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		eq	:	OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		q	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0);
		sclr	:	IN STD_LOGIC := '0';
		sload	:	IN STD_LOGIC := '0';
		sset	:	IN STD_LOGIC := '0';
		updown	:	IN STD_LOGIC := '1'
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_decode
	 GENERIC 
	 (
		LPM_DECODES	:	NATURAL;
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_decode"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		data	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		enable	:	IN STD_LOGIC := '1';
		eq	:	OUT STD_LOGIC_VECTOR(LPM_DECODES-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
 BEGIN

	wire_dprio_w_lg_w_lg_w_lg_s0_to_0694w695w696w(0) <= wire_dprio_w_lg_w_lg_s0_to_0694w695w(0) AND wire_state_mc_reg_w_q_range692w(0);
	wire_dprio_w_lg_w_lg_w_lg_s1_to_0713w714w715w(0) <= wire_dprio_w_lg_w_lg_s1_to_0713w714w(0) AND wire_state_mc_reg_w_q_range711w(0);
	wire_dprio_w_lg_w_lg_w_lg_s2_to_0729w730w731w(0) <= wire_dprio_w_lg_w_lg_s2_to_0729w730w(0) AND wire_state_mc_reg_w_q_range727w(0);
	wire_dprio_w_lg_w_lg_w_lg_wren683w706w719w(0) <= wire_dprio_w_lg_w_lg_wren683w706w(0) AND wire_dprio_w_lg_rdinc718w(0);
	wire_dprio_w_lg_w_lg_w_lg_wren683w706w707w(0) <= wire_dprio_w_lg_w_lg_wren683w706w(0) AND rden;
	wire_dprio_w_lg_w_lg_w_lg_wr_addr_state859w863w864w(0) <= wire_dprio_w_lg_w_lg_wr_addr_state859w863w(0) AND wire_pre_amble_cmpr_agb;
	wire_dprio_w_lg_w_lg_rd_data_output_state1039w1040w(0) <= wire_dprio_w_lg_rd_data_output_state1039w(0) AND wire_pre_amble_cmpr_agb;
	wire_dprio_w_lg_w_lg_wr_data_state974w975w(0) <= wire_dprio_w_lg_wr_data_state974w(0) AND wire_pre_amble_cmpr_agb;
	wire_dprio_w_lg_w_lg_s0_to_0694w695w(0) <= wire_dprio_w_lg_s0_to_0694w(0) AND wire_dprio_w_lg_s0_to_1693w(0);
	wire_dprio_w_lg_w_lg_s1_to_0713w714w(0) <= wire_dprio_w_lg_s1_to_0713w(0) AND wire_dprio_w_lg_s1_to_1712w(0);
	wire_dprio_w_lg_w_lg_s2_to_0729w730w(0) <= wire_dprio_w_lg_s2_to_0729w(0) AND wire_dprio_w_lg_s2_to_1728w(0);
	wire_dprio_w_lg_w_lg_wren683w706w(0) <= wire_dprio_w_lg_wren683w(0) AND wire_dprio_w_lg_wren_data705w(0);
	wire_dprio_w_lg_w_lg_wren683w684w(0) <= wire_dprio_w_lg_wren683w(0) AND wire_dprio_w_lg_w_lg_rden681w682w(0);
	wire_dprio_w_lg_w_lg_wren683w701w(0) <= wire_dprio_w_lg_wren683w(0) AND wire_dprio_w_lg_rdinc700w(0);
	wire_dprio_w_lg_w_lg_w_lg_w_lg_rden1095w1096w1097w1098w(0) <= wire_dprio_w_lg_w_lg_w_lg_rden1095w1096w1097w(0) AND wire_dprio_w_lg_startup_done1093w(0);
	wire_dprio_w_lg_w_lg_wr_addr_state859w863w(0) <= wire_dprio_w_lg_wr_addr_state859w(0) AND wire_addr_shift_reg_w_q_range862w(0);
	wire_dprio_w_lg_idle_state720w(0) <= idle_state AND wire_dprio_w_lg_w_lg_w_lg_wren683w706w719w(0);
	wire_dprio_w_lg_idle_state702w(0) <= idle_state AND wire_dprio_w_lg_w_lg_wren683w701w(0);
	wire_dprio_w_lg_idle_state709w(0) <= idle_state AND wire_dprio_w_lg_wren708w(0);
	wire_dprio_w_lg_idle_state686w(0) <= idle_state AND wire_dprio_w_lg_wren685w(0);
	wire_dprio_w_lg_idle_state723w(0) <= idle_state AND wire_dprio_w_lg_wren722w(0);
	wire_dprio_w_lg_rd_data_output_state1039w(0) <= rd_data_output_state AND wire_rd_out_data_shift_reg_w_q_range1038w(0);
	wire_dprio_w_lg_wr_data_state974w(0) <= wr_data_state AND wire_wr_out_data_shift_reg_w_q_range973w(0);
	wire_dprio_w_lg_s0_to_0694w(0) <= NOT s0_to_0;
	wire_dprio_w_lg_s0_to_1693w(0) <= NOT s0_to_1;
	wire_dprio_w_lg_s1_to_0713w(0) <= NOT s1_to_0;
	wire_dprio_w_lg_s1_to_1712w(0) <= NOT s1_to_1;
	wire_dprio_w_lg_s2_to_0729w(0) <= NOT s2_to_0;
	wire_dprio_w_lg_s2_to_1728w(0) <= NOT s2_to_1;
	wire_dprio_w_lg_startup_done1093w(0) <= NOT startup_done;
	wire_dprio_w_lg_startup_idle1094w(0) <= NOT startup_idle;
	wire_dprio_w_lg_wren683w(0) <= NOT wren;
	wire_dprio_w_lg_wren_data705w(0) <= NOT wren_data;
	wire_dprio_w_lg_w_lg_w_lg_rden1095w1096w1097w(0) <= wire_dprio_w_lg_w_lg_rden1095w1096w(0) OR wire_dprio_w_lg_startup_idle1094w(0);
	wire_dprio_w_lg_w_lg_rden681w682w(0) <= wire_dprio_w_lg_rden681w(0) OR wren_data;
	wire_dprio_w_lg_w_lg_rden1095w1096w(0) <= wire_dprio_w_lg_rden1095w(0) OR rdinc;
	wire_dprio_w_lg_rden681w(0) <= rden OR rdinc;
	wire_dprio_w_lg_rden1095w(0) <= rden OR wren;
	wire_dprio_w_lg_rdinc718w(0) <= rdinc OR rden;
	wire_dprio_w_lg_rdinc700w(0) <= rdinc OR wren_data;
	wire_dprio_w_lg_s0_to_1697w(0) <= s0_to_1 OR wire_dprio_w_lg_w_lg_w_lg_s0_to_0694w695w696w(0);
	wire_dprio_w_lg_s1_to_1716w(0) <= s1_to_1 OR wire_dprio_w_lg_w_lg_w_lg_s1_to_0713w714w715w(0);
	wire_dprio_w_lg_s2_to_1732w(0) <= s2_to_1 OR wire_dprio_w_lg_w_lg_w_lg_s2_to_0729w730w731w(0);
	wire_dprio_w_lg_wr_addr_state859w(0) <= wr_addr_state OR rd_addr_state;
	wire_dprio_w_lg_wren708w(0) <= wren OR wire_dprio_w_lg_w_lg_w_lg_wren683w706w707w(0);
	wire_dprio_w_lg_wren685w(0) <= wren OR wire_dprio_w_lg_w_lg_wren683w684w(0);
	wire_dprio_w_lg_wren722w(0) <= wren OR wren_data;
	busy <= busy_state;
	busy_state <= (write_state OR read_state);
	dataout <= in_data_shift_reg;
	dpriodisable <= (NOT wire_startup_cntr_w_lg_w_q_range1107w1116w(0));
	dprioin <= wire_dprioin_mux_dataout;
	dprioload <= (NOT (wire_startup_cntr_w_lg_w_q_range1099w1104w(0) AND (NOT startup_cntr(2))));
	idle_state <= wire_state_mc_decode_eq(0);
	rd_addr_done <= (rd_addr_state AND wire_state_mc_cmpr_aeb);
	rd_addr_state <= (wire_state_mc_decode_eq(5) AND startup_done);
	rd_data_done <= (rd_data_state AND wire_state_mc_cmpr_aeb);
	rd_data_input_state <= (wire_rd_data_output_cmpr_ageb AND rd_data_state);
	rd_data_output_state <= (wire_rd_data_output_cmpr_alb AND rd_data_state);
	rd_data_state <= (wire_state_mc_decode_eq(7) AND startup_done);
	rdinc <= '0';
	read_state <= (rd_addr_state OR rd_data_state);
	s0_to_0 <= ((wr_data_state AND wr_data_done) OR (rd_data_state AND rd_data_done));
	s0_to_1 <= ((wire_dprio_w_lg_idle_state686w(0) OR (wr_addr_state AND wr_addr_done)) OR (rd_addr_state AND rd_addr_done));
	s1_to_0 <= (((wr_data_state AND wr_data_done) OR (rd_data_state AND rd_data_done)) OR wire_dprio_w_lg_idle_state709w(0));
	s1_to_1 <= ((wire_dprio_w_lg_idle_state702w(0) OR (wr_addr_state AND wr_addr_done)) OR (rd_addr_state AND rd_addr_done));
	s2_to_0 <= ((((wr_addr_state AND wr_addr_done) OR (wr_data_state AND wr_data_done)) OR (rd_data_state AND rd_data_done)) OR wire_dprio_w_lg_idle_state723w(0));
	s2_to_1 <= (wire_dprio_w_lg_idle_state720w(0) OR (rd_addr_state AND rd_addr_done));
	startup_done <= (wire_startup_cntr_w_lg_w_q_range1107w1113w(0) AND startup_cntr(1));
	startup_idle <= (wire_startup_cntr_w_lg_w_q_range1099w1100w(0) AND (NOT (startup_cntr(2) XOR startup_cntr(1))));
	status_out <= ( rd_data_done & rd_addr_done & wr_data_done & wr_addr_done);
	wr_addr_done <= (wr_addr_state AND wire_state_mc_cmpr_aeb);
	wr_addr_state <= (wire_state_mc_decode_eq(1) AND startup_done);
	wr_data_done <= (wr_data_state AND wire_state_mc_cmpr_aeb);
	wr_data_state <= (wire_state_mc_decode_eq(3) AND startup_done);
	write_state <= (wr_addr_state OR wr_data_state);
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(0) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(0) <= wire_addr_shift_reg_asdata(0);
				ELSE addr_shift_reg(0) <= wire_addr_shift_reg_d(0);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(1) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(1) <= wire_addr_shift_reg_asdata(1);
				ELSE addr_shift_reg(1) <= wire_addr_shift_reg_d(1);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(2) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(2) <= wire_addr_shift_reg_asdata(2);
				ELSE addr_shift_reg(2) <= wire_addr_shift_reg_d(2);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(3) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(3) <= wire_addr_shift_reg_asdata(3);
				ELSE addr_shift_reg(3) <= wire_addr_shift_reg_d(3);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(4) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(4) <= wire_addr_shift_reg_asdata(4);
				ELSE addr_shift_reg(4) <= wire_addr_shift_reg_d(4);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(5) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(5) <= wire_addr_shift_reg_asdata(5);
				ELSE addr_shift_reg(5) <= wire_addr_shift_reg_d(5);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(6) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(6) <= wire_addr_shift_reg_asdata(6);
				ELSE addr_shift_reg(6) <= wire_addr_shift_reg_d(6);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(7) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(7) <= wire_addr_shift_reg_asdata(7);
				ELSE addr_shift_reg(7) <= wire_addr_shift_reg_d(7);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(8) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(8) <= wire_addr_shift_reg_asdata(8);
				ELSE addr_shift_reg(8) <= wire_addr_shift_reg_d(8);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(9) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(9) <= wire_addr_shift_reg_asdata(9);
				ELSE addr_shift_reg(9) <= wire_addr_shift_reg_d(9);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(10) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(10) <= wire_addr_shift_reg_asdata(10);
				ELSE addr_shift_reg(10) <= wire_addr_shift_reg_d(10);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(11) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(11) <= wire_addr_shift_reg_asdata(11);
				ELSE addr_shift_reg(11) <= wire_addr_shift_reg_d(11);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(12) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(12) <= wire_addr_shift_reg_asdata(12);
				ELSE addr_shift_reg(12) <= wire_addr_shift_reg_d(12);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(13) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(13) <= wire_addr_shift_reg_asdata(13);
				ELSE addr_shift_reg(13) <= wire_addr_shift_reg_d(13);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(14) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(14) <= wire_addr_shift_reg_asdata(14);
				ELSE addr_shift_reg(14) <= wire_addr_shift_reg_d(14);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(15) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(15) <= wire_addr_shift_reg_asdata(15);
				ELSE addr_shift_reg(15) <= wire_addr_shift_reg_d(15);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(16) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(16) <= wire_addr_shift_reg_asdata(16);
				ELSE addr_shift_reg(16) <= wire_addr_shift_reg_d(16);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(17) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(17) <= wire_addr_shift_reg_asdata(17);
				ELSE addr_shift_reg(17) <= wire_addr_shift_reg_d(17);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(18) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(18) <= wire_addr_shift_reg_asdata(18);
				ELSE addr_shift_reg(18) <= wire_addr_shift_reg_d(18);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(19) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(19) <= wire_addr_shift_reg_asdata(19);
				ELSE addr_shift_reg(19) <= wire_addr_shift_reg_d(19);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(20) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(20) <= wire_addr_shift_reg_asdata(20);
				ELSE addr_shift_reg(20) <= wire_addr_shift_reg_d(20);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(21) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(21) <= wire_addr_shift_reg_asdata(21);
				ELSE addr_shift_reg(21) <= wire_addr_shift_reg_d(21);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(22) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(22) <= wire_addr_shift_reg_asdata(22);
				ELSE addr_shift_reg(22) <= wire_addr_shift_reg_d(22);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(23) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(23) <= wire_addr_shift_reg_asdata(23);
				ELSE addr_shift_reg(23) <= wire_addr_shift_reg_d(23);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(24) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(24) <= wire_addr_shift_reg_asdata(24);
				ELSE addr_shift_reg(24) <= wire_addr_shift_reg_d(24);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(25) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(25) <= wire_addr_shift_reg_asdata(25);
				ELSE addr_shift_reg(25) <= wire_addr_shift_reg_d(25);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(26) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(26) <= wire_addr_shift_reg_asdata(26);
				ELSE addr_shift_reg(26) <= wire_addr_shift_reg_d(26);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(27) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(27) <= wire_addr_shift_reg_asdata(27);
				ELSE addr_shift_reg(27) <= wire_addr_shift_reg_d(27);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(28) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(28) <= wire_addr_shift_reg_asdata(28);
				ELSE addr_shift_reg(28) <= wire_addr_shift_reg_d(28);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(29) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(29) <= wire_addr_shift_reg_asdata(29);
				ELSE addr_shift_reg(29) <= wire_addr_shift_reg_d(29);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(30) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(30) <= wire_addr_shift_reg_asdata(30);
				ELSE addr_shift_reg(30) <= wire_addr_shift_reg_d(30);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(31) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(31) <= wire_addr_shift_reg_asdata(31);
				ELSE addr_shift_reg(31) <= wire_addr_shift_reg_d(31);
				END IF;
		END IF;
	END PROCESS;
	wire_addr_shift_reg_asdata <= ( "00" & "00" & "0" & quad_address(8 DOWNTO 0) & "10" & address);
	wire_addr_shift_reg_d <= ( addr_shift_reg(30 DOWNTO 0) & "0");
	wire_addr_shift_reg_w_q_range862w(0) <= addr_shift_reg(31);
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN in_data_shift_reg <= (OTHERS => '0');
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
			IF (rd_data_input_state = '1') THEN in_data_shift_reg <= ( in_data_shift_reg(14 DOWNTO 0) & dprioout);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(0) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(0) <= wire_rd_out_data_shift_reg_asdata(0);
				ELSE rd_out_data_shift_reg(0) <= wire_rd_out_data_shift_reg_d(0);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(1) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(1) <= wire_rd_out_data_shift_reg_asdata(1);
				ELSE rd_out_data_shift_reg(1) <= wire_rd_out_data_shift_reg_d(1);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(2) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(2) <= wire_rd_out_data_shift_reg_asdata(2);
				ELSE rd_out_data_shift_reg(2) <= wire_rd_out_data_shift_reg_d(2);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(3) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(3) <= wire_rd_out_data_shift_reg_asdata(3);
				ELSE rd_out_data_shift_reg(3) <= wire_rd_out_data_shift_reg_d(3);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(4) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(4) <= wire_rd_out_data_shift_reg_asdata(4);
				ELSE rd_out_data_shift_reg(4) <= wire_rd_out_data_shift_reg_d(4);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(5) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(5) <= wire_rd_out_data_shift_reg_asdata(5);
				ELSE rd_out_data_shift_reg(5) <= wire_rd_out_data_shift_reg_d(5);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(6) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(6) <= wire_rd_out_data_shift_reg_asdata(6);
				ELSE rd_out_data_shift_reg(6) <= wire_rd_out_data_shift_reg_d(6);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(7) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(7) <= wire_rd_out_data_shift_reg_asdata(7);
				ELSE rd_out_data_shift_reg(7) <= wire_rd_out_data_shift_reg_d(7);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(8) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(8) <= wire_rd_out_data_shift_reg_asdata(8);
				ELSE rd_out_data_shift_reg(8) <= wire_rd_out_data_shift_reg_d(8);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(9) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(9) <= wire_rd_out_data_shift_reg_asdata(9);
				ELSE rd_out_data_shift_reg(9) <= wire_rd_out_data_shift_reg_d(9);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(10) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(10) <= wire_rd_out_data_shift_reg_asdata(10);
				ELSE rd_out_data_shift_reg(10) <= wire_rd_out_data_shift_reg_d(10);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(11) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(11) <= wire_rd_out_data_shift_reg_asdata(11);
				ELSE rd_out_data_shift_reg(11) <= wire_rd_out_data_shift_reg_d(11);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(12) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(12) <= wire_rd_out_data_shift_reg_asdata(12);
				ELSE rd_out_data_shift_reg(12) <= wire_rd_out_data_shift_reg_d(12);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(13) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(13) <= wire_rd_out_data_shift_reg_asdata(13);
				ELSE rd_out_data_shift_reg(13) <= wire_rd_out_data_shift_reg_d(13);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(14) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(14) <= wire_rd_out_data_shift_reg_asdata(14);
				ELSE rd_out_data_shift_reg(14) <= wire_rd_out_data_shift_reg_d(14);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(15) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(15) <= wire_rd_out_data_shift_reg_asdata(15);
				ELSE rd_out_data_shift_reg(15) <= wire_rd_out_data_shift_reg_d(15);
				END IF;
		END IF;
	END PROCESS;
	wire_rd_out_data_shift_reg_asdata <= ( "00" & "1" & "1" & "0" & quad_address & "10");
	wire_rd_out_data_shift_reg_d <= ( rd_out_data_shift_reg(14 DOWNTO 0) & "0");
	wire_rd_out_data_shift_reg_w_q_range1038w(0) <= rd_out_data_shift_reg(15);
	PROCESS (dpclk)
	BEGIN
		IF (dpclk = '1' AND dpclk'event) THEN 
			IF (wire_startup_cntr_ena(0) = '1') THEN 
				IF (reset = '1') THEN startup_cntr(0) <= '0';
				ELSE startup_cntr(0) <= wire_startup_cntr_d(0);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk)
	BEGIN
		IF (dpclk = '1' AND dpclk'event) THEN 
			IF (wire_startup_cntr_ena(1) = '1') THEN 
				IF (reset = '1') THEN startup_cntr(1) <= '0';
				ELSE startup_cntr(1) <= wire_startup_cntr_d(1);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk)
	BEGIN
		IF (dpclk = '1' AND dpclk'event) THEN 
			IF (wire_startup_cntr_ena(2) = '1') THEN 
				IF (reset = '1') THEN startup_cntr(2) <= '0';
				ELSE startup_cntr(2) <= wire_startup_cntr_d(2);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	wire_startup_cntr_d <= ( wire_startup_cntr_w_lg_w_q_range1107w1108w & wire_startup_cntr_w_lg_w_q_range1099w1104w & wire_startup_cntr_w_lg_w_q_range1099w1100w);
	loop0 : FOR i IN 0 TO 2 GENERATE
		wire_startup_cntr_ena(i) <= wire_dprio_w_lg_w_lg_w_lg_w_lg_rden1095w1096w1097w1098w(0);
	END GENERATE loop0;
	wire_startup_cntr_w_lg_w_q_range1103w1106w(0) <= wire_startup_cntr_w_q_range1103w(0) AND wire_startup_cntr_w_q_range1099w(0);
	wire_startup_cntr_w_lg_w_q_range1107w1113w(0) <= wire_startup_cntr_w_q_range1107w(0) AND wire_startup_cntr_w_lg_w_q_range1099w1100w(0);
	wire_startup_cntr_w_lg_w_q_range1107w1116w(0) <= wire_startup_cntr_w_q_range1107w(0) AND wire_startup_cntr_w_lg_w_q_range1099w1115w(0);
	wire_startup_cntr_w_lg_w_q_range1099w1100w(0) <= NOT wire_startup_cntr_w_q_range1099w(0);
	wire_startup_cntr_w_lg_w_q_range1099w1115w(0) <= wire_startup_cntr_w_q_range1099w(0) OR wire_startup_cntr_w_q_range1103w(0);
	wire_startup_cntr_w_lg_w_q_range1099w1104w(0) <= wire_startup_cntr_w_q_range1099w(0) XOR wire_startup_cntr_w_q_range1103w(0);
	wire_startup_cntr_w_lg_w_q_range1107w1108w(0) <= wire_startup_cntr_w_q_range1107w(0) XOR wire_startup_cntr_w_lg_w_q_range1103w1106w(0);
	wire_startup_cntr_w_q_range1099w(0) <= startup_cntr(0);
	wire_startup_cntr_w_q_range1103w(0) <= startup_cntr(1);
	wire_startup_cntr_w_q_range1107w(0) <= startup_cntr(2);
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN state_mc_reg <= (OTHERS => '0');
		ELSIF (dpclk = '1' AND dpclk'event) THEN state_mc_reg <= ( wire_dprio_w_lg_s2_to_1732w & wire_dprio_w_lg_s1_to_1716w & wire_dprio_w_lg_s0_to_1697w);
		END IF;
	END PROCESS;
	wire_state_mc_reg_w_q_range692w(0) <= state_mc_reg(0);
	wire_state_mc_reg_w_q_range711w(0) <= state_mc_reg(1);
	wire_state_mc_reg_w_q_range727w(0) <= state_mc_reg(2);
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(0) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(0) <= wire_wr_out_data_shift_reg_asdata(0);
				ELSE wr_out_data_shift_reg(0) <= wire_wr_out_data_shift_reg_d(0);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(1) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(1) <= wire_wr_out_data_shift_reg_asdata(1);
				ELSE wr_out_data_shift_reg(1) <= wire_wr_out_data_shift_reg_d(1);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(2) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(2) <= wire_wr_out_data_shift_reg_asdata(2);
				ELSE wr_out_data_shift_reg(2) <= wire_wr_out_data_shift_reg_d(2);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(3) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(3) <= wire_wr_out_data_shift_reg_asdata(3);
				ELSE wr_out_data_shift_reg(3) <= wire_wr_out_data_shift_reg_d(3);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(4) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(4) <= wire_wr_out_data_shift_reg_asdata(4);
				ELSE wr_out_data_shift_reg(4) <= wire_wr_out_data_shift_reg_d(4);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(5) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(5) <= wire_wr_out_data_shift_reg_asdata(5);
				ELSE wr_out_data_shift_reg(5) <= wire_wr_out_data_shift_reg_d(5);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(6) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(6) <= wire_wr_out_data_shift_reg_asdata(6);
				ELSE wr_out_data_shift_reg(6) <= wire_wr_out_data_shift_reg_d(6);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(7) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(7) <= wire_wr_out_data_shift_reg_asdata(7);
				ELSE wr_out_data_shift_reg(7) <= wire_wr_out_data_shift_reg_d(7);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(8) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(8) <= wire_wr_out_data_shift_reg_asdata(8);
				ELSE wr_out_data_shift_reg(8) <= wire_wr_out_data_shift_reg_d(8);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(9) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(9) <= wire_wr_out_data_shift_reg_asdata(9);
				ELSE wr_out_data_shift_reg(9) <= wire_wr_out_data_shift_reg_d(9);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(10) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(10) <= wire_wr_out_data_shift_reg_asdata(10);
				ELSE wr_out_data_shift_reg(10) <= wire_wr_out_data_shift_reg_d(10);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(11) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(11) <= wire_wr_out_data_shift_reg_asdata(11);
				ELSE wr_out_data_shift_reg(11) <= wire_wr_out_data_shift_reg_d(11);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(12) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(12) <= wire_wr_out_data_shift_reg_asdata(12);
				ELSE wr_out_data_shift_reg(12) <= wire_wr_out_data_shift_reg_d(12);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(13) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(13) <= wire_wr_out_data_shift_reg_asdata(13);
				ELSE wr_out_data_shift_reg(13) <= wire_wr_out_data_shift_reg_d(13);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(14) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(14) <= wire_wr_out_data_shift_reg_asdata(14);
				ELSE wr_out_data_shift_reg(14) <= wire_wr_out_data_shift_reg_d(14);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(15) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(15) <= wire_wr_out_data_shift_reg_asdata(15);
				ELSE wr_out_data_shift_reg(15) <= wire_wr_out_data_shift_reg_d(15);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(16) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(16) <= wire_wr_out_data_shift_reg_asdata(16);
				ELSE wr_out_data_shift_reg(16) <= wire_wr_out_data_shift_reg_d(16);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(17) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(17) <= wire_wr_out_data_shift_reg_asdata(17);
				ELSE wr_out_data_shift_reg(17) <= wire_wr_out_data_shift_reg_d(17);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(18) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(18) <= wire_wr_out_data_shift_reg_asdata(18);
				ELSE wr_out_data_shift_reg(18) <= wire_wr_out_data_shift_reg_d(18);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(19) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(19) <= wire_wr_out_data_shift_reg_asdata(19);
				ELSE wr_out_data_shift_reg(19) <= wire_wr_out_data_shift_reg_d(19);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(20) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(20) <= wire_wr_out_data_shift_reg_asdata(20);
				ELSE wr_out_data_shift_reg(20) <= wire_wr_out_data_shift_reg_d(20);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(21) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(21) <= wire_wr_out_data_shift_reg_asdata(21);
				ELSE wr_out_data_shift_reg(21) <= wire_wr_out_data_shift_reg_d(21);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(22) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(22) <= wire_wr_out_data_shift_reg_asdata(22);
				ELSE wr_out_data_shift_reg(22) <= wire_wr_out_data_shift_reg_d(22);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(23) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(23) <= wire_wr_out_data_shift_reg_asdata(23);
				ELSE wr_out_data_shift_reg(23) <= wire_wr_out_data_shift_reg_d(23);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(24) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(24) <= wire_wr_out_data_shift_reg_asdata(24);
				ELSE wr_out_data_shift_reg(24) <= wire_wr_out_data_shift_reg_d(24);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(25) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(25) <= wire_wr_out_data_shift_reg_asdata(25);
				ELSE wr_out_data_shift_reg(25) <= wire_wr_out_data_shift_reg_d(25);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(26) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(26) <= wire_wr_out_data_shift_reg_asdata(26);
				ELSE wr_out_data_shift_reg(26) <= wire_wr_out_data_shift_reg_d(26);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(27) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(27) <= wire_wr_out_data_shift_reg_asdata(27);
				ELSE wr_out_data_shift_reg(27) <= wire_wr_out_data_shift_reg_d(27);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(28) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(28) <= wire_wr_out_data_shift_reg_asdata(28);
				ELSE wr_out_data_shift_reg(28) <= wire_wr_out_data_shift_reg_d(28);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(29) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(29) <= wire_wr_out_data_shift_reg_asdata(29);
				ELSE wr_out_data_shift_reg(29) <= wire_wr_out_data_shift_reg_d(29);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(30) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(30) <= wire_wr_out_data_shift_reg_asdata(30);
				ELSE wr_out_data_shift_reg(30) <= wire_wr_out_data_shift_reg_d(30);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(31) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(31) <= wire_wr_out_data_shift_reg_asdata(31);
				ELSE wr_out_data_shift_reg(31) <= wire_wr_out_data_shift_reg_d(31);
				END IF;
		END IF;
	END PROCESS;
	wire_wr_out_data_shift_reg_asdata <= ( "00" & "01" & "0" & quad_address(8 DOWNTO 0) & "10" & datain);
	wire_wr_out_data_shift_reg_d <= ( wr_out_data_shift_reg(30 DOWNTO 0) & "0");
	wire_wr_out_data_shift_reg_w_q_range973w(0) <= wr_out_data_shift_reg(31);
	wire_pre_amble_cmpr_w_lg_w_lg_agb860w1037w(0) <= wire_pre_amble_cmpr_w_lg_agb860w(0) AND rd_data_output_state;
	wire_pre_amble_cmpr_w_lg_w_lg_agb860w972w(0) <= wire_pre_amble_cmpr_w_lg_agb860w(0) AND wr_data_state;
	wire_pre_amble_cmpr_w_lg_agb860w(0) <= NOT wire_pre_amble_cmpr_agb;
	wire_pre_amble_cmpr_datab <= "011111";
	pre_amble_cmpr :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 6
	  )
	  PORT MAP ( 
		aeb => wire_pre_amble_cmpr_aeb,
		agb => wire_pre_amble_cmpr_agb,
		dataa => wire_state_mc_counter_q,
		datab => wire_pre_amble_cmpr_datab
	  );
	wire_rd_data_output_cmpr_datab <= "110000";
	rd_data_output_cmpr :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 6
	  )
	  PORT MAP ( 
		ageb => wire_rd_data_output_cmpr_ageb,
		alb => wire_rd_data_output_cmpr_alb,
		dataa => wire_state_mc_counter_q,
		datab => wire_rd_data_output_cmpr_datab
	  );
	wire_state_mc_cmpr_datab <= (OTHERS => '1');
	state_mc_cmpr :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 6
	  )
	  PORT MAP ( 
		aeb => wire_state_mc_cmpr_aeb,
		dataa => wire_state_mc_counter_q,
		datab => wire_state_mc_cmpr_datab
	  );
	wire_state_mc_counter_cnt_en <= wire_dprio_w_lg_write_state677w(0);
	wire_dprio_w_lg_write_state677w(0) <= write_state OR read_state;
	state_mc_counter :  lpm_counter
	  GENERIC MAP (
		lpm_port_updown => "PORT_UNUSED",
		lpm_width => 6
	  )
	  PORT MAP ( 
		clock => dpclk,
		cnt_en => wire_state_mc_counter_cnt_en,
		q => wire_state_mc_counter_q,
		sclr => reset
	  );
	state_mc_decode :  lpm_decode
	  GENERIC MAP (
		LPM_DECODES => 8,
		LPM_WIDTH => 3
	  )
	  PORT MAP ( 
		data => state_mc_reg,
		eq => wire_state_mc_decode_eq
	  );
	wire_dprioin_mux_dataout <= (((wire_dprio_w_lg_w_lg_w_lg_wr_addr_state859w863w864w(0) OR (wire_pre_amble_cmpr_w_lg_agb860w(0) AND wire_dprio_w_lg_wr_addr_state859w(0))) OR (wire_dprio_w_lg_w_lg_wr_data_state974w975w(0) OR wire_pre_amble_cmpr_w_lg_w_lg_agb860w972w(0))) OR (wire_dprio_w_lg_w_lg_rd_data_output_state1039w1040w(0) OR wire_pre_amble_cmpr_w_lg_w_lg_agb860w1037w(0))) OR NOT(((write_state OR rd_addr_state) OR rd_data_output_state));

 END RTL; --ALTGX_RECONFIG_CIV_alt_dprio_q9l


--lpm_mux CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone IV GX" LPM_SIZE=6 LPM_WIDTH=6 LPM_WIDTHS=3 data result sel
--VERSION_BEGIN 21.1 cbx_lpm_mux 2021:10:21:11:02:24:SJ cbx_mgl 2021:10:21:11:11:47:SJ  VERSION_END

--synthesis_resources = lut 30 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  ALTGX_RECONFIG_CIV_mux_cda IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (35 DOWNTO 0) := (OTHERS => '0');
		 result	:	OUT  STD_LOGIC_VECTOR (5 DOWNTO 0);
		 sel	:	IN  STD_LOGIC_VECTOR (2 DOWNTO 0) := (OTHERS => '0')
	 ); 
 END ALTGX_RECONFIG_CIV_mux_cda;

 ARCHITECTURE RTL OF ALTGX_RECONFIG_CIV_mux_cda IS

	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_lg_w_sel_node_range1128w1192w1193w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_lg_w_sel_node_range1128w1192w1261w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_lg_w_sel_node_range1128w1192w1328w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_lg_w_sel_node_range1128w1192w1395w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_lg_w_sel_node_range1128w1192w1462w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_lg_w_sel_node_range1128w1192w1529w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_result1155w1169w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_result1176w1186w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_result1224w1238w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_result1245w1255w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_result1291w1305w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_result1312w1322w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_result1358w1372w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_result1379w1389w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_result1425w1439w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_result1446w1456w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_result1492w1506w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_result1513w1523w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_sel_node_range1128w1194w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_sel_node_range1128w1262w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_sel_node_range1128w1329w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_sel_node_range1128w1396w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_sel_node_range1128w1463w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_sel_node_range1128w1530w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_data1149w_range1163w1164w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_data1150w_range1180w1181w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_data1218w_range1232w1233w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_data1219w_range1249w1250w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_data1285w_range1299w1300w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_data1286w_range1316w1317w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_data1352w_range1366w1367w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_data1353w_range1383w1384w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_data1419w_range1433w1434w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_data1420w_range1450w1451w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_data1486w_range1500w1501w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_data1487w_range1517w1518w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_sel1151w_range1159w1160w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_sel1151w_range1159w1179w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_sel1220w_range1228w1229w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_sel1220w_range1228w1248w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_sel1287w_range1295w1296w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_sel1287w_range1295w1315w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_sel1354w_range1362w1363w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_sel1354w_range1362w1382w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_sel1421w_range1429w1430w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_sel1421w_range1429w1449w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_sel1488w_range1496w1497w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_sel1488w_range1496w1516w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_result1155w1170w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_result1176w1187w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_result1224w1239w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_result1245w1256w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_result1291w1306w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_result1312w1323w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_result1358w1373w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_result1379w1390w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_result1425w1440w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_result1446w1457w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_result1492w1507w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_result1513w1524w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_sel_node_range1128w1192w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_sel1151w_range1157w1161w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_sel1151w_range1159w1162w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_sel1220w_range1226w1230w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_sel1220w_range1228w1231w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_sel1287w_range1293w1297w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_sel1287w_range1295w1298w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_sel1354w_range1360w1364w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_sel1354w_range1362w1365w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_sel1421w_range1427w1431w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_sel1421w_range1429w1432w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_sel1488w_range1494w1498w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_sel1488w_range1496w1499w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_data1149w_range1167w1168w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_data1150w_range1184w1185w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_data1218w_range1236w1237w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_data1219w_range1253w1254w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_data1285w_range1303w1304w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_data1286w_range1320w1321w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_data1352w_range1370w1371w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_data1353w_range1387w1388w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_data1419w_range1437w1438w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_data1420w_range1454w1455w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_data1486w_range1504w1505w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_data1487w_range1521w1522w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_sel1151w_range1157w1158w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_sel1151w_range1157w1178w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_sel1220w_range1226w1227w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_sel1220w_range1226w1247w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_sel1287w_range1293w1294w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_sel1287w_range1293w1314w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_sel1354w_range1360w1361w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_sel1354w_range1360w1381w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_sel1421w_range1427w1428w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_sel1421w_range1427w1448w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_sel1488w_range1494w1495w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_lg_w_w_sel1488w_range1494w1515w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  result_node :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  sel_ffs_wire :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  sel_node :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  w_data1129w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  w_data1149w :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  w_data1150w :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  w_data1198w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  w_data1218w :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  w_data1219w :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  w_data1265w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  w_data1285w :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  w_data1286w :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  w_data1332w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  w_data1352w :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  w_data1353w :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  w_data1399w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  w_data1419w :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  w_data1420w :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  w_data1466w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  w_data1486w :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  w_data1487w :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  w_result1130w :	STD_LOGIC;
	 SIGNAL  w_result1147w :	STD_LOGIC;
	 SIGNAL  w_result1148w :	STD_LOGIC;
	 SIGNAL  w_result1155w :	STD_LOGIC;
	 SIGNAL  w_result1176w :	STD_LOGIC;
	 SIGNAL  w_result1199w :	STD_LOGIC;
	 SIGNAL  w_result1216w :	STD_LOGIC;
	 SIGNAL  w_result1217w :	STD_LOGIC;
	 SIGNAL  w_result1224w :	STD_LOGIC;
	 SIGNAL  w_result1245w :	STD_LOGIC;
	 SIGNAL  w_result1266w :	STD_LOGIC;
	 SIGNAL  w_result1283w :	STD_LOGIC;
	 SIGNAL  w_result1284w :	STD_LOGIC;
	 SIGNAL  w_result1291w :	STD_LOGIC;
	 SIGNAL  w_result1312w :	STD_LOGIC;
	 SIGNAL  w_result1333w :	STD_LOGIC;
	 SIGNAL  w_result1350w :	STD_LOGIC;
	 SIGNAL  w_result1351w :	STD_LOGIC;
	 SIGNAL  w_result1358w :	STD_LOGIC;
	 SIGNAL  w_result1379w :	STD_LOGIC;
	 SIGNAL  w_result1400w :	STD_LOGIC;
	 SIGNAL  w_result1417w :	STD_LOGIC;
	 SIGNAL  w_result1418w :	STD_LOGIC;
	 SIGNAL  w_result1425w :	STD_LOGIC;
	 SIGNAL  w_result1446w :	STD_LOGIC;
	 SIGNAL  w_result1467w :	STD_LOGIC;
	 SIGNAL  w_result1484w :	STD_LOGIC;
	 SIGNAL  w_result1485w :	STD_LOGIC;
	 SIGNAL  w_result1492w :	STD_LOGIC;
	 SIGNAL  w_result1513w :	STD_LOGIC;
	 SIGNAL  w_sel1151w :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  w_sel1220w :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  w_sel1287w :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  w_sel1354w :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  w_sel1421w :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  w_sel1488w :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_sel_node_range1128w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_data1149w_range1163w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_data1149w_range1156w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_data1149w_range1167w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_data1150w_range1180w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_data1150w_range1177w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_data1150w_range1184w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_data1218w_range1232w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_data1218w_range1225w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_data1218w_range1236w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_data1219w_range1249w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_data1219w_range1246w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_data1219w_range1253w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_data1285w_range1299w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_data1285w_range1292w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_data1285w_range1303w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_data1286w_range1316w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_data1286w_range1313w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_data1286w_range1320w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_data1352w_range1366w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_data1352w_range1359w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_data1352w_range1370w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_data1353w_range1383w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_data1353w_range1380w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_data1353w_range1387w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_data1419w_range1433w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_data1419w_range1426w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_data1419w_range1437w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_data1420w_range1450w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_data1420w_range1447w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_data1420w_range1454w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_data1486w_range1500w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_data1486w_range1493w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_data1486w_range1504w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_data1487w_range1517w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_data1487w_range1514w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_data1487w_range1521w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_sel1151w_range1157w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_sel1151w_range1159w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_sel1220w_range1226w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_sel1220w_range1228w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_sel1287w_range1293w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_sel1287w_range1295w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_sel1354w_range1360w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_sel1354w_range1362w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_sel1421w_range1427w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_sel1421w_range1429w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_sel1488w_range1494w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_w_w_sel1488w_range1496w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
 BEGIN

	wire_central_pcs_first_word_mux_w_lg_w_lg_w_sel_node_range1128w1192w1193w(0) <= wire_central_pcs_first_word_mux_w_lg_w_sel_node_range1128w1192w(0) AND w_result1147w;
	wire_central_pcs_first_word_mux_w_lg_w_lg_w_sel_node_range1128w1192w1261w(0) <= wire_central_pcs_first_word_mux_w_lg_w_sel_node_range1128w1192w(0) AND w_result1216w;
	wire_central_pcs_first_word_mux_w_lg_w_lg_w_sel_node_range1128w1192w1328w(0) <= wire_central_pcs_first_word_mux_w_lg_w_sel_node_range1128w1192w(0) AND w_result1283w;
	wire_central_pcs_first_word_mux_w_lg_w_lg_w_sel_node_range1128w1192w1395w(0) <= wire_central_pcs_first_word_mux_w_lg_w_sel_node_range1128w1192w(0) AND w_result1350w;
	wire_central_pcs_first_word_mux_w_lg_w_lg_w_sel_node_range1128w1192w1462w(0) <= wire_central_pcs_first_word_mux_w_lg_w_sel_node_range1128w1192w(0) AND w_result1417w;
	wire_central_pcs_first_word_mux_w_lg_w_lg_w_sel_node_range1128w1192w1529w(0) <= wire_central_pcs_first_word_mux_w_lg_w_sel_node_range1128w1192w(0) AND w_result1484w;
	wire_central_pcs_first_word_mux_w_lg_w_result1155w1169w(0) <= w_result1155w AND wire_central_pcs_first_word_mux_w_lg_w_w_data1149w_range1167w1168w(0);
	wire_central_pcs_first_word_mux_w_lg_w_result1176w1186w(0) <= w_result1176w AND wire_central_pcs_first_word_mux_w_lg_w_w_data1150w_range1184w1185w(0);
	wire_central_pcs_first_word_mux_w_lg_w_result1224w1238w(0) <= w_result1224w AND wire_central_pcs_first_word_mux_w_lg_w_w_data1218w_range1236w1237w(0);
	wire_central_pcs_first_word_mux_w_lg_w_result1245w1255w(0) <= w_result1245w AND wire_central_pcs_first_word_mux_w_lg_w_w_data1219w_range1253w1254w(0);
	wire_central_pcs_first_word_mux_w_lg_w_result1291w1305w(0) <= w_result1291w AND wire_central_pcs_first_word_mux_w_lg_w_w_data1285w_range1303w1304w(0);
	wire_central_pcs_first_word_mux_w_lg_w_result1312w1322w(0) <= w_result1312w AND wire_central_pcs_first_word_mux_w_lg_w_w_data1286w_range1320w1321w(0);
	wire_central_pcs_first_word_mux_w_lg_w_result1358w1372w(0) <= w_result1358w AND wire_central_pcs_first_word_mux_w_lg_w_w_data1352w_range1370w1371w(0);
	wire_central_pcs_first_word_mux_w_lg_w_result1379w1389w(0) <= w_result1379w AND wire_central_pcs_first_word_mux_w_lg_w_w_data1353w_range1387w1388w(0);
	wire_central_pcs_first_word_mux_w_lg_w_result1425w1439w(0) <= w_result1425w AND wire_central_pcs_first_word_mux_w_lg_w_w_data1419w_range1437w1438w(0);
	wire_central_pcs_first_word_mux_w_lg_w_result1446w1456w(0) <= w_result1446w AND wire_central_pcs_first_word_mux_w_lg_w_w_data1420w_range1454w1455w(0);
	wire_central_pcs_first_word_mux_w_lg_w_result1492w1506w(0) <= w_result1492w AND wire_central_pcs_first_word_mux_w_lg_w_w_data1486w_range1504w1505w(0);
	wire_central_pcs_first_word_mux_w_lg_w_result1513w1523w(0) <= w_result1513w AND wire_central_pcs_first_word_mux_w_lg_w_w_data1487w_range1521w1522w(0);
	wire_central_pcs_first_word_mux_w_lg_w_sel_node_range1128w1194w(0) <= wire_central_pcs_first_word_mux_w_sel_node_range1128w(0) AND w_result1148w;
	wire_central_pcs_first_word_mux_w_lg_w_sel_node_range1128w1262w(0) <= wire_central_pcs_first_word_mux_w_sel_node_range1128w(0) AND w_result1217w;
	wire_central_pcs_first_word_mux_w_lg_w_sel_node_range1128w1329w(0) <= wire_central_pcs_first_word_mux_w_sel_node_range1128w(0) AND w_result1284w;
	wire_central_pcs_first_word_mux_w_lg_w_sel_node_range1128w1396w(0) <= wire_central_pcs_first_word_mux_w_sel_node_range1128w(0) AND w_result1351w;
	wire_central_pcs_first_word_mux_w_lg_w_sel_node_range1128w1463w(0) <= wire_central_pcs_first_word_mux_w_sel_node_range1128w(0) AND w_result1418w;
	wire_central_pcs_first_word_mux_w_lg_w_sel_node_range1128w1530w(0) <= wire_central_pcs_first_word_mux_w_sel_node_range1128w(0) AND w_result1485w;
	wire_central_pcs_first_word_mux_w_lg_w_w_data1149w_range1163w1164w(0) <= wire_central_pcs_first_word_mux_w_w_data1149w_range1163w(0) AND wire_central_pcs_first_word_mux_w_lg_w_w_sel1151w_range1159w1162w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_data1150w_range1180w1181w(0) <= wire_central_pcs_first_word_mux_w_w_data1150w_range1180w(0) AND wire_central_pcs_first_word_mux_w_lg_w_w_sel1151w_range1159w1162w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_data1218w_range1232w1233w(0) <= wire_central_pcs_first_word_mux_w_w_data1218w_range1232w(0) AND wire_central_pcs_first_word_mux_w_lg_w_w_sel1220w_range1228w1231w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_data1219w_range1249w1250w(0) <= wire_central_pcs_first_word_mux_w_w_data1219w_range1249w(0) AND wire_central_pcs_first_word_mux_w_lg_w_w_sel1220w_range1228w1231w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_data1285w_range1299w1300w(0) <= wire_central_pcs_first_word_mux_w_w_data1285w_range1299w(0) AND wire_central_pcs_first_word_mux_w_lg_w_w_sel1287w_range1295w1298w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_data1286w_range1316w1317w(0) <= wire_central_pcs_first_word_mux_w_w_data1286w_range1316w(0) AND wire_central_pcs_first_word_mux_w_lg_w_w_sel1287w_range1295w1298w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_data1352w_range1366w1367w(0) <= wire_central_pcs_first_word_mux_w_w_data1352w_range1366w(0) AND wire_central_pcs_first_word_mux_w_lg_w_w_sel1354w_range1362w1365w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_data1353w_range1383w1384w(0) <= wire_central_pcs_first_word_mux_w_w_data1353w_range1383w(0) AND wire_central_pcs_first_word_mux_w_lg_w_w_sel1354w_range1362w1365w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_data1419w_range1433w1434w(0) <= wire_central_pcs_first_word_mux_w_w_data1419w_range1433w(0) AND wire_central_pcs_first_word_mux_w_lg_w_w_sel1421w_range1429w1432w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_data1420w_range1450w1451w(0) <= wire_central_pcs_first_word_mux_w_w_data1420w_range1450w(0) AND wire_central_pcs_first_word_mux_w_lg_w_w_sel1421w_range1429w1432w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_data1486w_range1500w1501w(0) <= wire_central_pcs_first_word_mux_w_w_data1486w_range1500w(0) AND wire_central_pcs_first_word_mux_w_lg_w_w_sel1488w_range1496w1499w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_data1487w_range1517w1518w(0) <= wire_central_pcs_first_word_mux_w_w_data1487w_range1517w(0) AND wire_central_pcs_first_word_mux_w_lg_w_w_sel1488w_range1496w1499w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_sel1151w_range1159w1160w(0) <= wire_central_pcs_first_word_mux_w_w_sel1151w_range1159w(0) AND wire_central_pcs_first_word_mux_w_lg_w_w_sel1151w_range1157w1158w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_sel1151w_range1159w1179w(0) <= wire_central_pcs_first_word_mux_w_w_sel1151w_range1159w(0) AND wire_central_pcs_first_word_mux_w_lg_w_w_sel1151w_range1157w1178w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_sel1220w_range1228w1229w(0) <= wire_central_pcs_first_word_mux_w_w_sel1220w_range1228w(0) AND wire_central_pcs_first_word_mux_w_lg_w_w_sel1220w_range1226w1227w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_sel1220w_range1228w1248w(0) <= wire_central_pcs_first_word_mux_w_w_sel1220w_range1228w(0) AND wire_central_pcs_first_word_mux_w_lg_w_w_sel1220w_range1226w1247w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_sel1287w_range1295w1296w(0) <= wire_central_pcs_first_word_mux_w_w_sel1287w_range1295w(0) AND wire_central_pcs_first_word_mux_w_lg_w_w_sel1287w_range1293w1294w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_sel1287w_range1295w1315w(0) <= wire_central_pcs_first_word_mux_w_w_sel1287w_range1295w(0) AND wire_central_pcs_first_word_mux_w_lg_w_w_sel1287w_range1293w1314w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_sel1354w_range1362w1363w(0) <= wire_central_pcs_first_word_mux_w_w_sel1354w_range1362w(0) AND wire_central_pcs_first_word_mux_w_lg_w_w_sel1354w_range1360w1361w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_sel1354w_range1362w1382w(0) <= wire_central_pcs_first_word_mux_w_w_sel1354w_range1362w(0) AND wire_central_pcs_first_word_mux_w_lg_w_w_sel1354w_range1360w1381w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_sel1421w_range1429w1430w(0) <= wire_central_pcs_first_word_mux_w_w_sel1421w_range1429w(0) AND wire_central_pcs_first_word_mux_w_lg_w_w_sel1421w_range1427w1428w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_sel1421w_range1429w1449w(0) <= wire_central_pcs_first_word_mux_w_w_sel1421w_range1429w(0) AND wire_central_pcs_first_word_mux_w_lg_w_w_sel1421w_range1427w1448w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_sel1488w_range1496w1497w(0) <= wire_central_pcs_first_word_mux_w_w_sel1488w_range1496w(0) AND wire_central_pcs_first_word_mux_w_lg_w_w_sel1488w_range1494w1495w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_sel1488w_range1496w1516w(0) <= wire_central_pcs_first_word_mux_w_w_sel1488w_range1496w(0) AND wire_central_pcs_first_word_mux_w_lg_w_w_sel1488w_range1494w1515w(0);
	wire_central_pcs_first_word_mux_w_lg_w_result1155w1170w(0) <= NOT w_result1155w;
	wire_central_pcs_first_word_mux_w_lg_w_result1176w1187w(0) <= NOT w_result1176w;
	wire_central_pcs_first_word_mux_w_lg_w_result1224w1239w(0) <= NOT w_result1224w;
	wire_central_pcs_first_word_mux_w_lg_w_result1245w1256w(0) <= NOT w_result1245w;
	wire_central_pcs_first_word_mux_w_lg_w_result1291w1306w(0) <= NOT w_result1291w;
	wire_central_pcs_first_word_mux_w_lg_w_result1312w1323w(0) <= NOT w_result1312w;
	wire_central_pcs_first_word_mux_w_lg_w_result1358w1373w(0) <= NOT w_result1358w;
	wire_central_pcs_first_word_mux_w_lg_w_result1379w1390w(0) <= NOT w_result1379w;
	wire_central_pcs_first_word_mux_w_lg_w_result1425w1440w(0) <= NOT w_result1425w;
	wire_central_pcs_first_word_mux_w_lg_w_result1446w1457w(0) <= NOT w_result1446w;
	wire_central_pcs_first_word_mux_w_lg_w_result1492w1507w(0) <= NOT w_result1492w;
	wire_central_pcs_first_word_mux_w_lg_w_result1513w1524w(0) <= NOT w_result1513w;
	wire_central_pcs_first_word_mux_w_lg_w_sel_node_range1128w1192w(0) <= NOT wire_central_pcs_first_word_mux_w_sel_node_range1128w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_sel1151w_range1157w1161w(0) <= NOT wire_central_pcs_first_word_mux_w_w_sel1151w_range1157w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_sel1151w_range1159w1162w(0) <= NOT wire_central_pcs_first_word_mux_w_w_sel1151w_range1159w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_sel1220w_range1226w1230w(0) <= NOT wire_central_pcs_first_word_mux_w_w_sel1220w_range1226w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_sel1220w_range1228w1231w(0) <= NOT wire_central_pcs_first_word_mux_w_w_sel1220w_range1228w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_sel1287w_range1293w1297w(0) <= NOT wire_central_pcs_first_word_mux_w_w_sel1287w_range1293w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_sel1287w_range1295w1298w(0) <= NOT wire_central_pcs_first_word_mux_w_w_sel1287w_range1295w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_sel1354w_range1360w1364w(0) <= NOT wire_central_pcs_first_word_mux_w_w_sel1354w_range1360w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_sel1354w_range1362w1365w(0) <= NOT wire_central_pcs_first_word_mux_w_w_sel1354w_range1362w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_sel1421w_range1427w1431w(0) <= NOT wire_central_pcs_first_word_mux_w_w_sel1421w_range1427w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_sel1421w_range1429w1432w(0) <= NOT wire_central_pcs_first_word_mux_w_w_sel1421w_range1429w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_sel1488w_range1494w1498w(0) <= NOT wire_central_pcs_first_word_mux_w_w_sel1488w_range1494w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_sel1488w_range1496w1499w(0) <= NOT wire_central_pcs_first_word_mux_w_w_sel1488w_range1496w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_data1149w_range1167w1168w(0) <= wire_central_pcs_first_word_mux_w_w_data1149w_range1167w(0) OR wire_central_pcs_first_word_mux_w_lg_w_w_sel1151w_range1157w1161w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_data1150w_range1184w1185w(0) <= wire_central_pcs_first_word_mux_w_w_data1150w_range1184w(0) OR wire_central_pcs_first_word_mux_w_lg_w_w_sel1151w_range1157w1161w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_data1218w_range1236w1237w(0) <= wire_central_pcs_first_word_mux_w_w_data1218w_range1236w(0) OR wire_central_pcs_first_word_mux_w_lg_w_w_sel1220w_range1226w1230w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_data1219w_range1253w1254w(0) <= wire_central_pcs_first_word_mux_w_w_data1219w_range1253w(0) OR wire_central_pcs_first_word_mux_w_lg_w_w_sel1220w_range1226w1230w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_data1285w_range1303w1304w(0) <= wire_central_pcs_first_word_mux_w_w_data1285w_range1303w(0) OR wire_central_pcs_first_word_mux_w_lg_w_w_sel1287w_range1293w1297w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_data1286w_range1320w1321w(0) <= wire_central_pcs_first_word_mux_w_w_data1286w_range1320w(0) OR wire_central_pcs_first_word_mux_w_lg_w_w_sel1287w_range1293w1297w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_data1352w_range1370w1371w(0) <= wire_central_pcs_first_word_mux_w_w_data1352w_range1370w(0) OR wire_central_pcs_first_word_mux_w_lg_w_w_sel1354w_range1360w1364w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_data1353w_range1387w1388w(0) <= wire_central_pcs_first_word_mux_w_w_data1353w_range1387w(0) OR wire_central_pcs_first_word_mux_w_lg_w_w_sel1354w_range1360w1364w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_data1419w_range1437w1438w(0) <= wire_central_pcs_first_word_mux_w_w_data1419w_range1437w(0) OR wire_central_pcs_first_word_mux_w_lg_w_w_sel1421w_range1427w1431w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_data1420w_range1454w1455w(0) <= wire_central_pcs_first_word_mux_w_w_data1420w_range1454w(0) OR wire_central_pcs_first_word_mux_w_lg_w_w_sel1421w_range1427w1431w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_data1486w_range1504w1505w(0) <= wire_central_pcs_first_word_mux_w_w_data1486w_range1504w(0) OR wire_central_pcs_first_word_mux_w_lg_w_w_sel1488w_range1494w1498w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_data1487w_range1521w1522w(0) <= wire_central_pcs_first_word_mux_w_w_data1487w_range1521w(0) OR wire_central_pcs_first_word_mux_w_lg_w_w_sel1488w_range1494w1498w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_sel1151w_range1157w1158w(0) <= wire_central_pcs_first_word_mux_w_w_sel1151w_range1157w(0) OR wire_central_pcs_first_word_mux_w_w_data1149w_range1156w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_sel1151w_range1157w1178w(0) <= wire_central_pcs_first_word_mux_w_w_sel1151w_range1157w(0) OR wire_central_pcs_first_word_mux_w_w_data1150w_range1177w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_sel1220w_range1226w1227w(0) <= wire_central_pcs_first_word_mux_w_w_sel1220w_range1226w(0) OR wire_central_pcs_first_word_mux_w_w_data1218w_range1225w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_sel1220w_range1226w1247w(0) <= wire_central_pcs_first_word_mux_w_w_sel1220w_range1226w(0) OR wire_central_pcs_first_word_mux_w_w_data1219w_range1246w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_sel1287w_range1293w1294w(0) <= wire_central_pcs_first_word_mux_w_w_sel1287w_range1293w(0) OR wire_central_pcs_first_word_mux_w_w_data1285w_range1292w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_sel1287w_range1293w1314w(0) <= wire_central_pcs_first_word_mux_w_w_sel1287w_range1293w(0) OR wire_central_pcs_first_word_mux_w_w_data1286w_range1313w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_sel1354w_range1360w1361w(0) <= wire_central_pcs_first_word_mux_w_w_sel1354w_range1360w(0) OR wire_central_pcs_first_word_mux_w_w_data1352w_range1359w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_sel1354w_range1360w1381w(0) <= wire_central_pcs_first_word_mux_w_w_sel1354w_range1360w(0) OR wire_central_pcs_first_word_mux_w_w_data1353w_range1380w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_sel1421w_range1427w1428w(0) <= wire_central_pcs_first_word_mux_w_w_sel1421w_range1427w(0) OR wire_central_pcs_first_word_mux_w_w_data1419w_range1426w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_sel1421w_range1427w1448w(0) <= wire_central_pcs_first_word_mux_w_w_sel1421w_range1427w(0) OR wire_central_pcs_first_word_mux_w_w_data1420w_range1447w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_sel1488w_range1494w1495w(0) <= wire_central_pcs_first_word_mux_w_w_sel1488w_range1494w(0) OR wire_central_pcs_first_word_mux_w_w_data1486w_range1493w(0);
	wire_central_pcs_first_word_mux_w_lg_w_w_sel1488w_range1494w1515w(0) <= wire_central_pcs_first_word_mux_w_w_sel1488w_range1494w(0) OR wire_central_pcs_first_word_mux_w_w_data1487w_range1514w(0);
	result <= result_node;
	result_node <= ( w_result1467w & w_result1400w & w_result1333w & w_result1266w & w_result1199w & w_result1130w);
	sel_ffs_wire <= ( sel(2 DOWNTO 0));
	sel_node <= ( sel_ffs_wire(2) & sel(1 DOWNTO 0));
	w_data1129w <= ( "00" & data(30) & data(24) & data(18) & data(12) & data(6) & data(0));
	w_data1149w <= w_data1129w(3 DOWNTO 0);
	w_data1150w <= w_data1129w(7 DOWNTO 4);
	w_data1198w <= ( "00" & data(31) & data(25) & data(19) & data(13) & data(7) & data(1));
	w_data1218w <= w_data1198w(3 DOWNTO 0);
	w_data1219w <= w_data1198w(7 DOWNTO 4);
	w_data1265w <= ( "00" & data(32) & data(26) & data(20) & data(14) & data(8) & data(2));
	w_data1285w <= w_data1265w(3 DOWNTO 0);
	w_data1286w <= w_data1265w(7 DOWNTO 4);
	w_data1332w <= ( "00" & data(33) & data(27) & data(21) & data(15) & data(9) & data(3));
	w_data1352w <= w_data1332w(3 DOWNTO 0);
	w_data1353w <= w_data1332w(7 DOWNTO 4);
	w_data1399w <= ( "00" & data(34) & data(28) & data(22) & data(16) & data(10) & data(4));
	w_data1419w <= w_data1399w(3 DOWNTO 0);
	w_data1420w <= w_data1399w(7 DOWNTO 4);
	w_data1466w <= ( "00" & data(35) & data(29) & data(23) & data(17) & data(11) & data(5));
	w_data1486w <= w_data1466w(3 DOWNTO 0);
	w_data1487w <= w_data1466w(7 DOWNTO 4);
	w_result1130w <= (wire_central_pcs_first_word_mux_w_lg_w_sel_node_range1128w1194w(0) OR wire_central_pcs_first_word_mux_w_lg_w_lg_w_sel_node_range1128w1192w1193w(0));
	w_result1147w <= (((w_data1149w(1) AND w_sel1151w(0)) AND wire_central_pcs_first_word_mux_w_lg_w_result1155w1170w(0)) OR wire_central_pcs_first_word_mux_w_lg_w_result1155w1169w(0));
	w_result1148w <= (((w_data1150w(1) AND w_sel1151w(0)) AND wire_central_pcs_first_word_mux_w_lg_w_result1176w1187w(0)) OR wire_central_pcs_first_word_mux_w_lg_w_result1176w1186w(0));
	w_result1155w <= ((wire_central_pcs_first_word_mux_w_lg_w_w_data1149w_range1163w1164w(0) AND wire_central_pcs_first_word_mux_w_lg_w_w_sel1151w_range1157w1161w(0)) OR wire_central_pcs_first_word_mux_w_lg_w_w_sel1151w_range1159w1160w(0));
	w_result1176w <= ((wire_central_pcs_first_word_mux_w_lg_w_w_data1150w_range1180w1181w(0) AND wire_central_pcs_first_word_mux_w_lg_w_w_sel1151w_range1157w1161w(0)) OR wire_central_pcs_first_word_mux_w_lg_w_w_sel1151w_range1159w1179w(0));
	w_result1199w <= (wire_central_pcs_first_word_mux_w_lg_w_sel_node_range1128w1262w(0) OR wire_central_pcs_first_word_mux_w_lg_w_lg_w_sel_node_range1128w1192w1261w(0));
	w_result1216w <= (((w_data1218w(1) AND w_sel1220w(0)) AND wire_central_pcs_first_word_mux_w_lg_w_result1224w1239w(0)) OR wire_central_pcs_first_word_mux_w_lg_w_result1224w1238w(0));
	w_result1217w <= (((w_data1219w(1) AND w_sel1220w(0)) AND wire_central_pcs_first_word_mux_w_lg_w_result1245w1256w(0)) OR wire_central_pcs_first_word_mux_w_lg_w_result1245w1255w(0));
	w_result1224w <= ((wire_central_pcs_first_word_mux_w_lg_w_w_data1218w_range1232w1233w(0) AND wire_central_pcs_first_word_mux_w_lg_w_w_sel1220w_range1226w1230w(0)) OR wire_central_pcs_first_word_mux_w_lg_w_w_sel1220w_range1228w1229w(0));
	w_result1245w <= ((wire_central_pcs_first_word_mux_w_lg_w_w_data1219w_range1249w1250w(0) AND wire_central_pcs_first_word_mux_w_lg_w_w_sel1220w_range1226w1230w(0)) OR wire_central_pcs_first_word_mux_w_lg_w_w_sel1220w_range1228w1248w(0));
	w_result1266w <= (wire_central_pcs_first_word_mux_w_lg_w_sel_node_range1128w1329w(0) OR wire_central_pcs_first_word_mux_w_lg_w_lg_w_sel_node_range1128w1192w1328w(0));
	w_result1283w <= (((w_data1285w(1) AND w_sel1287w(0)) AND wire_central_pcs_first_word_mux_w_lg_w_result1291w1306w(0)) OR wire_central_pcs_first_word_mux_w_lg_w_result1291w1305w(0));
	w_result1284w <= (((w_data1286w(1) AND w_sel1287w(0)) AND wire_central_pcs_first_word_mux_w_lg_w_result1312w1323w(0)) OR wire_central_pcs_first_word_mux_w_lg_w_result1312w1322w(0));
	w_result1291w <= ((wire_central_pcs_first_word_mux_w_lg_w_w_data1285w_range1299w1300w(0) AND wire_central_pcs_first_word_mux_w_lg_w_w_sel1287w_range1293w1297w(0)) OR wire_central_pcs_first_word_mux_w_lg_w_w_sel1287w_range1295w1296w(0));
	w_result1312w <= ((wire_central_pcs_first_word_mux_w_lg_w_w_data1286w_range1316w1317w(0) AND wire_central_pcs_first_word_mux_w_lg_w_w_sel1287w_range1293w1297w(0)) OR wire_central_pcs_first_word_mux_w_lg_w_w_sel1287w_range1295w1315w(0));
	w_result1333w <= (wire_central_pcs_first_word_mux_w_lg_w_sel_node_range1128w1396w(0) OR wire_central_pcs_first_word_mux_w_lg_w_lg_w_sel_node_range1128w1192w1395w(0));
	w_result1350w <= (((w_data1352w(1) AND w_sel1354w(0)) AND wire_central_pcs_first_word_mux_w_lg_w_result1358w1373w(0)) OR wire_central_pcs_first_word_mux_w_lg_w_result1358w1372w(0));
	w_result1351w <= (((w_data1353w(1) AND w_sel1354w(0)) AND wire_central_pcs_first_word_mux_w_lg_w_result1379w1390w(0)) OR wire_central_pcs_first_word_mux_w_lg_w_result1379w1389w(0));
	w_result1358w <= ((wire_central_pcs_first_word_mux_w_lg_w_w_data1352w_range1366w1367w(0) AND wire_central_pcs_first_word_mux_w_lg_w_w_sel1354w_range1360w1364w(0)) OR wire_central_pcs_first_word_mux_w_lg_w_w_sel1354w_range1362w1363w(0));
	w_result1379w <= ((wire_central_pcs_first_word_mux_w_lg_w_w_data1353w_range1383w1384w(0) AND wire_central_pcs_first_word_mux_w_lg_w_w_sel1354w_range1360w1364w(0)) OR wire_central_pcs_first_word_mux_w_lg_w_w_sel1354w_range1362w1382w(0));
	w_result1400w <= (wire_central_pcs_first_word_mux_w_lg_w_sel_node_range1128w1463w(0) OR wire_central_pcs_first_word_mux_w_lg_w_lg_w_sel_node_range1128w1192w1462w(0));
	w_result1417w <= (((w_data1419w(1) AND w_sel1421w(0)) AND wire_central_pcs_first_word_mux_w_lg_w_result1425w1440w(0)) OR wire_central_pcs_first_word_mux_w_lg_w_result1425w1439w(0));
	w_result1418w <= (((w_data1420w(1) AND w_sel1421w(0)) AND wire_central_pcs_first_word_mux_w_lg_w_result1446w1457w(0)) OR wire_central_pcs_first_word_mux_w_lg_w_result1446w1456w(0));
	w_result1425w <= ((wire_central_pcs_first_word_mux_w_lg_w_w_data1419w_range1433w1434w(0) AND wire_central_pcs_first_word_mux_w_lg_w_w_sel1421w_range1427w1431w(0)) OR wire_central_pcs_first_word_mux_w_lg_w_w_sel1421w_range1429w1430w(0));
	w_result1446w <= ((wire_central_pcs_first_word_mux_w_lg_w_w_data1420w_range1450w1451w(0) AND wire_central_pcs_first_word_mux_w_lg_w_w_sel1421w_range1427w1431w(0)) OR wire_central_pcs_first_word_mux_w_lg_w_w_sel1421w_range1429w1449w(0));
	w_result1467w <= (wire_central_pcs_first_word_mux_w_lg_w_sel_node_range1128w1530w(0) OR wire_central_pcs_first_word_mux_w_lg_w_lg_w_sel_node_range1128w1192w1529w(0));
	w_result1484w <= (((w_data1486w(1) AND w_sel1488w(0)) AND wire_central_pcs_first_word_mux_w_lg_w_result1492w1507w(0)) OR wire_central_pcs_first_word_mux_w_lg_w_result1492w1506w(0));
	w_result1485w <= (((w_data1487w(1) AND w_sel1488w(0)) AND wire_central_pcs_first_word_mux_w_lg_w_result1513w1524w(0)) OR wire_central_pcs_first_word_mux_w_lg_w_result1513w1523w(0));
	w_result1492w <= ((wire_central_pcs_first_word_mux_w_lg_w_w_data1486w_range1500w1501w(0) AND wire_central_pcs_first_word_mux_w_lg_w_w_sel1488w_range1494w1498w(0)) OR wire_central_pcs_first_word_mux_w_lg_w_w_sel1488w_range1496w1497w(0));
	w_result1513w <= ((wire_central_pcs_first_word_mux_w_lg_w_w_data1487w_range1517w1518w(0) AND wire_central_pcs_first_word_mux_w_lg_w_w_sel1488w_range1494w1498w(0)) OR wire_central_pcs_first_word_mux_w_lg_w_w_sel1488w_range1496w1516w(0));
	w_sel1151w <= sel_node(1 DOWNTO 0);
	w_sel1220w <= sel_node(1 DOWNTO 0);
	w_sel1287w <= sel_node(1 DOWNTO 0);
	w_sel1354w <= sel_node(1 DOWNTO 0);
	w_sel1421w <= sel_node(1 DOWNTO 0);
	w_sel1488w <= sel_node(1 DOWNTO 0);
	wire_central_pcs_first_word_mux_w_sel_node_range1128w(0) <= sel_node(2);
	wire_central_pcs_first_word_mux_w_w_data1149w_range1163w(0) <= w_data1149w(0);
	wire_central_pcs_first_word_mux_w_w_data1149w_range1156w(0) <= w_data1149w(2);
	wire_central_pcs_first_word_mux_w_w_data1149w_range1167w(0) <= w_data1149w(3);
	wire_central_pcs_first_word_mux_w_w_data1150w_range1180w(0) <= w_data1150w(0);
	wire_central_pcs_first_word_mux_w_w_data1150w_range1177w(0) <= w_data1150w(2);
	wire_central_pcs_first_word_mux_w_w_data1150w_range1184w(0) <= w_data1150w(3);
	wire_central_pcs_first_word_mux_w_w_data1218w_range1232w(0) <= w_data1218w(0);
	wire_central_pcs_first_word_mux_w_w_data1218w_range1225w(0) <= w_data1218w(2);
	wire_central_pcs_first_word_mux_w_w_data1218w_range1236w(0) <= w_data1218w(3);
	wire_central_pcs_first_word_mux_w_w_data1219w_range1249w(0) <= w_data1219w(0);
	wire_central_pcs_first_word_mux_w_w_data1219w_range1246w(0) <= w_data1219w(2);
	wire_central_pcs_first_word_mux_w_w_data1219w_range1253w(0) <= w_data1219w(3);
	wire_central_pcs_first_word_mux_w_w_data1285w_range1299w(0) <= w_data1285w(0);
	wire_central_pcs_first_word_mux_w_w_data1285w_range1292w(0) <= w_data1285w(2);
	wire_central_pcs_first_word_mux_w_w_data1285w_range1303w(0) <= w_data1285w(3);
	wire_central_pcs_first_word_mux_w_w_data1286w_range1316w(0) <= w_data1286w(0);
	wire_central_pcs_first_word_mux_w_w_data1286w_range1313w(0) <= w_data1286w(2);
	wire_central_pcs_first_word_mux_w_w_data1286w_range1320w(0) <= w_data1286w(3);
	wire_central_pcs_first_word_mux_w_w_data1352w_range1366w(0) <= w_data1352w(0);
	wire_central_pcs_first_word_mux_w_w_data1352w_range1359w(0) <= w_data1352w(2);
	wire_central_pcs_first_word_mux_w_w_data1352w_range1370w(0) <= w_data1352w(3);
	wire_central_pcs_first_word_mux_w_w_data1353w_range1383w(0) <= w_data1353w(0);
	wire_central_pcs_first_word_mux_w_w_data1353w_range1380w(0) <= w_data1353w(2);
	wire_central_pcs_first_word_mux_w_w_data1353w_range1387w(0) <= w_data1353w(3);
	wire_central_pcs_first_word_mux_w_w_data1419w_range1433w(0) <= w_data1419w(0);
	wire_central_pcs_first_word_mux_w_w_data1419w_range1426w(0) <= w_data1419w(2);
	wire_central_pcs_first_word_mux_w_w_data1419w_range1437w(0) <= w_data1419w(3);
	wire_central_pcs_first_word_mux_w_w_data1420w_range1450w(0) <= w_data1420w(0);
	wire_central_pcs_first_word_mux_w_w_data1420w_range1447w(0) <= w_data1420w(2);
	wire_central_pcs_first_word_mux_w_w_data1420w_range1454w(0) <= w_data1420w(3);
	wire_central_pcs_first_word_mux_w_w_data1486w_range1500w(0) <= w_data1486w(0);
	wire_central_pcs_first_word_mux_w_w_data1486w_range1493w(0) <= w_data1486w(2);
	wire_central_pcs_first_word_mux_w_w_data1486w_range1504w(0) <= w_data1486w(3);
	wire_central_pcs_first_word_mux_w_w_data1487w_range1517w(0) <= w_data1487w(0);
	wire_central_pcs_first_word_mux_w_w_data1487w_range1514w(0) <= w_data1487w(2);
	wire_central_pcs_first_word_mux_w_w_data1487w_range1521w(0) <= w_data1487w(3);
	wire_central_pcs_first_word_mux_w_w_sel1151w_range1157w(0) <= w_sel1151w(0);
	wire_central_pcs_first_word_mux_w_w_sel1151w_range1159w(0) <= w_sel1151w(1);
	wire_central_pcs_first_word_mux_w_w_sel1220w_range1226w(0) <= w_sel1220w(0);
	wire_central_pcs_first_word_mux_w_w_sel1220w_range1228w(0) <= w_sel1220w(1);
	wire_central_pcs_first_word_mux_w_w_sel1287w_range1293w(0) <= w_sel1287w(0);
	wire_central_pcs_first_word_mux_w_w_sel1287w_range1295w(0) <= w_sel1287w(1);
	wire_central_pcs_first_word_mux_w_w_sel1354w_range1360w(0) <= w_sel1354w(0);
	wire_central_pcs_first_word_mux_w_w_sel1354w_range1362w(0) <= w_sel1354w(1);
	wire_central_pcs_first_word_mux_w_w_sel1421w_range1427w(0) <= w_sel1421w(0);
	wire_central_pcs_first_word_mux_w_w_sel1421w_range1429w(0) <= w_sel1421w(1);
	wire_central_pcs_first_word_mux_w_w_sel1488w_range1494w(0) <= w_sel1488w(0);
	wire_central_pcs_first_word_mux_w_w_sel1488w_range1496w(0) <= w_sel1488w(1);

 END RTL; --ALTGX_RECONFIG_CIV_mux_cda


--lpm_mux CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone IV GX" LPM_SIZE=4 LPM_WIDTH=5 LPM_WIDTHS=2 data result sel
--VERSION_BEGIN 21.1 cbx_lpm_mux 2021:10:21:11:02:24:SJ cbx_mgl 2021:10:21:11:11:47:SJ  VERSION_END

--synthesis_resources = lut 10 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  ALTGX_RECONFIG_CIV_mux_8da IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (19 DOWNTO 0) := (OTHERS => '0');
		 result	:	OUT  STD_LOGIC_VECTOR (4 DOWNTO 0);
		 sel	:	IN  STD_LOGIC_VECTOR (1 DOWNTO 0) := (OTHERS => '0')
	 ); 
 END ALTGX_RECONFIG_CIV_mux_8da;

 ARCHITECTURE RTL OF ALTGX_RECONFIG_CIV_mux_8da IS

	 SIGNAL  wire_max_word_per_mif_type_w_lg_w_result1548w1559w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_lg_w_result1578w1585w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_lg_w_result1603w1610w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_lg_w_result1628w1635w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_lg_w_result1653w1660w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_lg_w_sel_node_range1551w1552w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_lg_w_sel_node_range1551w1580w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_lg_w_sel_node_range1551w1605w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_lg_w_sel_node_range1551w1630w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_lg_w_sel_node_range1551w1655w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_lg_w_w_data1536w_range1539w1555w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_lg_w_w_data1566w_range1569w1581w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_lg_w_w_data1591w_range1594w1606w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_lg_w_w_data1616w_range1619w1631w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_lg_w_w_data1641w_range1644w1656w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_lg_w_result1548w1560w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_lg_w_result1578w1586w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_lg_w_result1603w1611w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_lg_w_result1628w1636w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_lg_w_result1653w1661w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_lg_w_sel_node_range1549w1553w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_lg_w_sel_node_range1551w1554w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_lg_w_sel_node_range1549w1550w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_lg_w_sel_node_range1549w1579w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_lg_w_sel_node_range1549w1604w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_lg_w_sel_node_range1549w1629w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_lg_w_sel_node_range1549w1654w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_lg_w_w_data1536w_range1546w1558w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_lg_w_w_data1566w_range1576w1584w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_lg_w_w_data1591w_range1601w1609w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_lg_w_w_data1616w_range1626w1634w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_lg_w_w_data1641w_range1651w1659w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  result_node :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  sel_node :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  w_data1536w :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  w_data1566w :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  w_data1591w :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  w_data1616w :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  w_data1641w :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  w_result1537w :	STD_LOGIC;
	 SIGNAL  w_result1548w :	STD_LOGIC;
	 SIGNAL  w_result1567w :	STD_LOGIC;
	 SIGNAL  w_result1578w :	STD_LOGIC;
	 SIGNAL  w_result1592w :	STD_LOGIC;
	 SIGNAL  w_result1603w :	STD_LOGIC;
	 SIGNAL  w_result1617w :	STD_LOGIC;
	 SIGNAL  w_result1628w :	STD_LOGIC;
	 SIGNAL  w_result1642w :	STD_LOGIC;
	 SIGNAL  w_result1653w :	STD_LOGIC;
	 SIGNAL  wire_max_word_per_mif_type_w_sel_node_range1549w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_sel_node_range1551w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_w_data1536w_range1539w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_w_data1536w_range1544w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_w_data1536w_range1546w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_w_data1566w_range1569w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_w_data1566w_range1574w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_w_data1566w_range1576w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_w_data1591w_range1594w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_w_data1591w_range1599w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_w_data1591w_range1601w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_w_data1616w_range1619w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_w_data1616w_range1624w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_w_data1616w_range1626w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_w_data1641w_range1644w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_w_data1641w_range1649w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_w_w_data1641w_range1651w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
 BEGIN

	wire_max_word_per_mif_type_w_lg_w_result1548w1559w(0) <= w_result1548w AND wire_max_word_per_mif_type_w_lg_w_w_data1536w_range1546w1558w(0);
	wire_max_word_per_mif_type_w_lg_w_result1578w1585w(0) <= w_result1578w AND wire_max_word_per_mif_type_w_lg_w_w_data1566w_range1576w1584w(0);
	wire_max_word_per_mif_type_w_lg_w_result1603w1610w(0) <= w_result1603w AND wire_max_word_per_mif_type_w_lg_w_w_data1591w_range1601w1609w(0);
	wire_max_word_per_mif_type_w_lg_w_result1628w1635w(0) <= w_result1628w AND wire_max_word_per_mif_type_w_lg_w_w_data1616w_range1626w1634w(0);
	wire_max_word_per_mif_type_w_lg_w_result1653w1660w(0) <= w_result1653w AND wire_max_word_per_mif_type_w_lg_w_w_data1641w_range1651w1659w(0);
	wire_max_word_per_mif_type_w_lg_w_sel_node_range1551w1552w(0) <= wire_max_word_per_mif_type_w_sel_node_range1551w(0) AND wire_max_word_per_mif_type_w_lg_w_sel_node_range1549w1550w(0);
	wire_max_word_per_mif_type_w_lg_w_sel_node_range1551w1580w(0) <= wire_max_word_per_mif_type_w_sel_node_range1551w(0) AND wire_max_word_per_mif_type_w_lg_w_sel_node_range1549w1579w(0);
	wire_max_word_per_mif_type_w_lg_w_sel_node_range1551w1605w(0) <= wire_max_word_per_mif_type_w_sel_node_range1551w(0) AND wire_max_word_per_mif_type_w_lg_w_sel_node_range1549w1604w(0);
	wire_max_word_per_mif_type_w_lg_w_sel_node_range1551w1630w(0) <= wire_max_word_per_mif_type_w_sel_node_range1551w(0) AND wire_max_word_per_mif_type_w_lg_w_sel_node_range1549w1629w(0);
	wire_max_word_per_mif_type_w_lg_w_sel_node_range1551w1655w(0) <= wire_max_word_per_mif_type_w_sel_node_range1551w(0) AND wire_max_word_per_mif_type_w_lg_w_sel_node_range1549w1654w(0);
	wire_max_word_per_mif_type_w_lg_w_w_data1536w_range1539w1555w(0) <= wire_max_word_per_mif_type_w_w_data1536w_range1539w(0) AND wire_max_word_per_mif_type_w_lg_w_sel_node_range1551w1554w(0);
	wire_max_word_per_mif_type_w_lg_w_w_data1566w_range1569w1581w(0) <= wire_max_word_per_mif_type_w_w_data1566w_range1569w(0) AND wire_max_word_per_mif_type_w_lg_w_sel_node_range1551w1554w(0);
	wire_max_word_per_mif_type_w_lg_w_w_data1591w_range1594w1606w(0) <= wire_max_word_per_mif_type_w_w_data1591w_range1594w(0) AND wire_max_word_per_mif_type_w_lg_w_sel_node_range1551w1554w(0);
	wire_max_word_per_mif_type_w_lg_w_w_data1616w_range1619w1631w(0) <= wire_max_word_per_mif_type_w_w_data1616w_range1619w(0) AND wire_max_word_per_mif_type_w_lg_w_sel_node_range1551w1554w(0);
	wire_max_word_per_mif_type_w_lg_w_w_data1641w_range1644w1656w(0) <= wire_max_word_per_mif_type_w_w_data1641w_range1644w(0) AND wire_max_word_per_mif_type_w_lg_w_sel_node_range1551w1554w(0);
	wire_max_word_per_mif_type_w_lg_w_result1548w1560w(0) <= NOT w_result1548w;
	wire_max_word_per_mif_type_w_lg_w_result1578w1586w(0) <= NOT w_result1578w;
	wire_max_word_per_mif_type_w_lg_w_result1603w1611w(0) <= NOT w_result1603w;
	wire_max_word_per_mif_type_w_lg_w_result1628w1636w(0) <= NOT w_result1628w;
	wire_max_word_per_mif_type_w_lg_w_result1653w1661w(0) <= NOT w_result1653w;
	wire_max_word_per_mif_type_w_lg_w_sel_node_range1549w1553w(0) <= NOT wire_max_word_per_mif_type_w_sel_node_range1549w(0);
	wire_max_word_per_mif_type_w_lg_w_sel_node_range1551w1554w(0) <= NOT wire_max_word_per_mif_type_w_sel_node_range1551w(0);
	wire_max_word_per_mif_type_w_lg_w_sel_node_range1549w1550w(0) <= wire_max_word_per_mif_type_w_sel_node_range1549w(0) OR wire_max_word_per_mif_type_w_w_data1536w_range1544w(0);
	wire_max_word_per_mif_type_w_lg_w_sel_node_range1549w1579w(0) <= wire_max_word_per_mif_type_w_sel_node_range1549w(0) OR wire_max_word_per_mif_type_w_w_data1566w_range1574w(0);
	wire_max_word_per_mif_type_w_lg_w_sel_node_range1549w1604w(0) <= wire_max_word_per_mif_type_w_sel_node_range1549w(0) OR wire_max_word_per_mif_type_w_w_data1591w_range1599w(0);
	wire_max_word_per_mif_type_w_lg_w_sel_node_range1549w1629w(0) <= wire_max_word_per_mif_type_w_sel_node_range1549w(0) OR wire_max_word_per_mif_type_w_w_data1616w_range1624w(0);
	wire_max_word_per_mif_type_w_lg_w_sel_node_range1549w1654w(0) <= wire_max_word_per_mif_type_w_sel_node_range1549w(0) OR wire_max_word_per_mif_type_w_w_data1641w_range1649w(0);
	wire_max_word_per_mif_type_w_lg_w_w_data1536w_range1546w1558w(0) <= wire_max_word_per_mif_type_w_w_data1536w_range1546w(0) OR wire_max_word_per_mif_type_w_lg_w_sel_node_range1549w1553w(0);
	wire_max_word_per_mif_type_w_lg_w_w_data1566w_range1576w1584w(0) <= wire_max_word_per_mif_type_w_w_data1566w_range1576w(0) OR wire_max_word_per_mif_type_w_lg_w_sel_node_range1549w1553w(0);
	wire_max_word_per_mif_type_w_lg_w_w_data1591w_range1601w1609w(0) <= wire_max_word_per_mif_type_w_w_data1591w_range1601w(0) OR wire_max_word_per_mif_type_w_lg_w_sel_node_range1549w1553w(0);
	wire_max_word_per_mif_type_w_lg_w_w_data1616w_range1626w1634w(0) <= wire_max_word_per_mif_type_w_w_data1616w_range1626w(0) OR wire_max_word_per_mif_type_w_lg_w_sel_node_range1549w1553w(0);
	wire_max_word_per_mif_type_w_lg_w_w_data1641w_range1651w1659w(0) <= wire_max_word_per_mif_type_w_w_data1641w_range1651w(0) OR wire_max_word_per_mif_type_w_lg_w_sel_node_range1549w1553w(0);
	result <= result_node;
	result_node <= ( w_result1642w & w_result1617w & w_result1592w & w_result1567w & w_result1537w);
	sel_node <= ( sel(1 DOWNTO 0));
	w_data1536w <= ( data(15) & data(10) & data(5) & data(0));
	w_data1566w <= ( data(16) & data(11) & data(6) & data(1));
	w_data1591w <= ( data(17) & data(12) & data(7) & data(2));
	w_data1616w <= ( data(18) & data(13) & data(8) & data(3));
	w_data1641w <= ( data(19) & data(14) & data(9) & data(4));
	w_result1537w <= (((w_data1536w(1) AND sel_node(0)) AND wire_max_word_per_mif_type_w_lg_w_result1548w1560w(0)) OR wire_max_word_per_mif_type_w_lg_w_result1548w1559w(0));
	w_result1548w <= ((wire_max_word_per_mif_type_w_lg_w_w_data1536w_range1539w1555w(0) AND wire_max_word_per_mif_type_w_lg_w_sel_node_range1549w1553w(0)) OR wire_max_word_per_mif_type_w_lg_w_sel_node_range1551w1552w(0));
	w_result1567w <= (((w_data1566w(1) AND sel_node(0)) AND wire_max_word_per_mif_type_w_lg_w_result1578w1586w(0)) OR wire_max_word_per_mif_type_w_lg_w_result1578w1585w(0));
	w_result1578w <= ((wire_max_word_per_mif_type_w_lg_w_w_data1566w_range1569w1581w(0) AND wire_max_word_per_mif_type_w_lg_w_sel_node_range1549w1553w(0)) OR wire_max_word_per_mif_type_w_lg_w_sel_node_range1551w1580w(0));
	w_result1592w <= (((w_data1591w(1) AND sel_node(0)) AND wire_max_word_per_mif_type_w_lg_w_result1603w1611w(0)) OR wire_max_word_per_mif_type_w_lg_w_result1603w1610w(0));
	w_result1603w <= ((wire_max_word_per_mif_type_w_lg_w_w_data1591w_range1594w1606w(0) AND wire_max_word_per_mif_type_w_lg_w_sel_node_range1549w1553w(0)) OR wire_max_word_per_mif_type_w_lg_w_sel_node_range1551w1605w(0));
	w_result1617w <= (((w_data1616w(1) AND sel_node(0)) AND wire_max_word_per_mif_type_w_lg_w_result1628w1636w(0)) OR wire_max_word_per_mif_type_w_lg_w_result1628w1635w(0));
	w_result1628w <= ((wire_max_word_per_mif_type_w_lg_w_w_data1616w_range1619w1631w(0) AND wire_max_word_per_mif_type_w_lg_w_sel_node_range1549w1553w(0)) OR wire_max_word_per_mif_type_w_lg_w_sel_node_range1551w1630w(0));
	w_result1642w <= (((w_data1641w(1) AND sel_node(0)) AND wire_max_word_per_mif_type_w_lg_w_result1653w1661w(0)) OR wire_max_word_per_mif_type_w_lg_w_result1653w1660w(0));
	w_result1653w <= ((wire_max_word_per_mif_type_w_lg_w_w_data1641w_range1644w1656w(0) AND wire_max_word_per_mif_type_w_lg_w_sel_node_range1549w1553w(0)) OR wire_max_word_per_mif_type_w_lg_w_sel_node_range1551w1655w(0));
	wire_max_word_per_mif_type_w_sel_node_range1549w(0) <= sel_node(0);
	wire_max_word_per_mif_type_w_sel_node_range1551w(0) <= sel_node(1);
	wire_max_word_per_mif_type_w_w_data1536w_range1539w(0) <= w_data1536w(0);
	wire_max_word_per_mif_type_w_w_data1536w_range1544w(0) <= w_data1536w(2);
	wire_max_word_per_mif_type_w_w_data1536w_range1546w(0) <= w_data1536w(3);
	wire_max_word_per_mif_type_w_w_data1566w_range1569w(0) <= w_data1566w(0);
	wire_max_word_per_mif_type_w_w_data1566w_range1574w(0) <= w_data1566w(2);
	wire_max_word_per_mif_type_w_w_data1566w_range1576w(0) <= w_data1566w(3);
	wire_max_word_per_mif_type_w_w_data1591w_range1594w(0) <= w_data1591w(0);
	wire_max_word_per_mif_type_w_w_data1591w_range1599w(0) <= w_data1591w(2);
	wire_max_word_per_mif_type_w_w_data1591w_range1601w(0) <= w_data1591w(3);
	wire_max_word_per_mif_type_w_w_data1616w_range1619w(0) <= w_data1616w(0);
	wire_max_word_per_mif_type_w_w_data1616w_range1624w(0) <= w_data1616w(2);
	wire_max_word_per_mif_type_w_w_data1616w_range1626w(0) <= w_data1616w(3);
	wire_max_word_per_mif_type_w_w_data1641w_range1644w(0) <= w_data1641w(0);
	wire_max_word_per_mif_type_w_w_data1641w_range1649w(0) <= w_data1641w(2);
	wire_max_word_per_mif_type_w_w_data1641w_range1651w(0) <= w_data1641w(3);

 END RTL; --ALTGX_RECONFIG_CIV_mux_8da

 LIBRARY altera_mf;
 USE altera_mf.all;

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = alt_cal_c3gxb 1 lpm_add_sub 1 lpm_compare 22 lpm_counter 4 lpm_decode 2 lut 41 reg 166 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  ALTGX_RECONFIG_CIV_alt_c3gxb_reconfig_osa1 IS 
	 PORT 
	 ( 
		 busy	:	OUT  STD_LOGIC;
		 channel_reconfig_done	:	OUT  STD_LOGIC;
		 error	:	OUT  STD_LOGIC;
		 reconfig_address_en	:	OUT  STD_LOGIC;
		 reconfig_address_out	:	OUT  STD_LOGIC_VECTOR (5 DOWNTO 0);
		 reconfig_clk	:	IN  STD_LOGIC;
		 reconfig_data	:	IN  STD_LOGIC_VECTOR (15 DOWNTO 0) := (OTHERS => '0');
		 reconfig_fromgxb	:	IN  STD_LOGIC_VECTOR (4 DOWNTO 0);
		 reconfig_mode_sel	:	IN  STD_LOGIC_VECTOR (2 DOWNTO 0) := (OTHERS => '0');
		 reconfig_reset	:	IN  STD_LOGIC := '0';
		 reconfig_togxb	:	OUT  STD_LOGIC_VECTOR (3 DOWNTO 0);
		 write_all	:	IN  STD_LOGIC := '0'
	 ); 
 END ALTGX_RECONFIG_CIV_alt_c3gxb_reconfig_osa1;

 ARCHITECTURE RTL OF ALTGX_RECONFIG_CIV_alt_c3gxb_reconfig_osa1 IS

	 ATTRIBUTE synthesis_clearbox : natural;
	 ATTRIBUTE synthesis_clearbox OF RTL : ARCHITECTURE IS 2;
	 ATTRIBUTE ALTERA_ATTRIBUTE : string;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF RTL : ARCHITECTURE IS "{-to address_pres_reg[11]} DPRIO_CHANNEL_NUM=11;{-to address_pres_reg[10]} DPRIO_CHANNEL_NUM=10;{-to address_pres_reg[9]} DPRIO_CHANNEL_NUM=9;{-to address_pres_reg[8]} DPRIO_CHANNEL_NUM=8;{-to address_pres_reg[7]} DPRIO_CHANNEL_NUM=7;{-to address_pres_reg[6]} DPRIO_CHANNEL_NUM=6;{-to address_pres_reg[5]} DPRIO_CHANNEL_NUM=5;{-to address_pres_reg[4]} DPRIO_CHANNEL_NUM=4;{-to address_pres_reg[3]} DPRIO_CHANNEL_NUM=3;{-to address_pres_reg[2]} DPRIO_CHANNEL_NUM=2;{-to address_pres_reg[1]} DPRIO_CHANNEL_NUM=1;{-to address_pres_reg[0]} DPRIO_CHANNEL_NUM=0";

	 SIGNAL  wire_calibration_c3gxb_w_lg_w_lg_busy97w101w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_calibration_c3gxb_w_lg_w_lg_busy97w98w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_calibration_c3gxb_w_lg_w_lg_busy97w104w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_calibration_c3gxb_w_lg_w_lg_busy97w107w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_calibration_c3gxb_w_lg_w_lg_busy97w110w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_calibration_c3gxb_w_lg_busy102w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_calibration_c3gxb_w_lg_busy99w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_calibration_c3gxb_w_lg_busy97w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_calibration_c3gxb_busy	:	STD_LOGIC;
	 SIGNAL  wire_calibration_c3gxb_dprio_addr	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_calibration_c3gxb_dprio_dataout	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_calibration_c3gxb_dprio_rden	:	STD_LOGIC;
	 SIGNAL  wire_calibration_c3gxb_dprio_wren	:	STD_LOGIC;
	 SIGNAL  wire_calibration_c3gxb_quad_addr	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_calibration_c3gxb_reset	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_offset_cancellation_reset82w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_calibration_c3gxb_retain_addr	:	STD_LOGIC;
	 SIGNAL  wire_dprio_w_lg_w_lg_w_status_out_range382w404w405w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_busy125w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_status_out_range382w404w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_address	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_calibration_c3gxb_w_lg_w_lg_busy102w103w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_dprio_busy	:	STD_LOGIC;
	 SIGNAL  wire_dprio_datain	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_calibration_c3gxb_w_lg_w_lg_busy99w100w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_dprio_dataout	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_dprio_dpriodisable	:	STD_LOGIC;
	 SIGNAL  wire_dprio_dprioin	:	STD_LOGIC;
	 SIGNAL  wire_dprio_dprioload	:	STD_LOGIC;
	 SIGNAL  wire_dprio_rden	:	STD_LOGIC;
	 SIGNAL  wire_calibration_c3gxb_w_lg_w_lg_busy105w106w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_status_out	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_dprio_wren	:	STD_LOGIC;
	 SIGNAL  wire_calibration_c3gxb_w_lg_w_lg_busy108w109w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_wren_data	:	STD_LOGIC;
	 SIGNAL  wire_calibration_c3gxb_w_lg_w_lg_busy111w112w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_status_out_range382w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_status_out_range403w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 address_pres_reg	:	STD_LOGIC_VECTOR(11 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF address_pres_reg : SIGNAL IS "PRESERVE_REGISTER=ON";

	 SIGNAL  wire_address_pres_reg_w_lg_w_lg_w_q_range66w67w68w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_address_pres_reg_w_lg_w_q_range70w71w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_address_pres_reg_w_lg_w_q_range66w67w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_address_pres_reg_w_lg_w_lg_w_lg_w_q_range66w67w68w69w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_address_pres_reg_w_q_range64w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_address_pres_reg_w_q_range70w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_address_pres_reg_w_q_range65w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_address_pres_reg_w_q_range66w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 delay_mif_head	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF delay_mif_head : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL	 wire_delay_mif_head_ena	:	STD_LOGIC;
	 SIGNAL	 delay_second_mif_head	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF delay_second_mif_head : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL	 wire_delay_second_mif_head_ena	:	STD_LOGIC;
	 SIGNAL	 dprio_dataout_reg	:	STD_LOGIC_VECTOR(15 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF dprio_dataout_reg : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL  wire_dprio_dataout_reg_w_q_range226w	:	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  wire_dprio_dataout_reg_w_q_range264w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_dprio_dataout_reg_w_q_range251w	:	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  wire_dprio_dataout_reg_w_q_range218w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_dprio_dataout_reg_w_q_range234w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_dprio_dataout_reg_w_q_range288w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_dprio_dataout_reg_w_q_range257w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_dprio_dataout_reg_w_q_range209w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_dataout_reg_w_q_range267w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_dprio_dataout_reg_w_q_range242w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_dprio_dataout_reg_w_q_range312w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_dprio_dataout_reg_w_q_range276w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_dprio_dataout_reg_w_q_range297w	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_dprio_dataout_reg_w_q_range321w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 dprio_pulse_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF dprio_pulse_reg : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL	 wire_dprio_pulse_reg_ena	:	STD_LOGIC;
	 SIGNAL	 end_mif_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF end_mif_reg : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL	 error_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 is_illegal_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 mif_central_pcs_error_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF mif_central_pcs_error_reg : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL	 wire_mif_central_pcs_error_reg_clrn	:	STD_LOGIC;
	 SIGNAL	 mif_stage	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF mif_stage : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL	 wire_mif_stage_sclr	:	STD_LOGIC;
	 SIGNAL  wire_mif_stage_w_lg_q194w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 wire_mif_type_reg_d	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL	 mif_type_reg	:	STD_LOGIC_VECTOR(3 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF mif_type_reg : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL	 wire_mif_type_reg_ena	:	STD_LOGIC_VECTOR(3 DOWNTO 0);
	 SIGNAL	 wire_mif_type_reg_sclr	:	STD_LOGIC_VECTOR(3 DOWNTO 0);
	 SIGNAL  wire_mif_type_reg_w_lg_w575w576w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_mif_type_reg_w_lg_w_lg_w_lg_w_lg_w_q_range492w571w572w573w574w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_mif_type_reg_w_lg_w_q_range504w505w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_mif_type_reg_w_lg_w_q_range499w500w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_mif_type_reg_w_lg_w_q_range495w496w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_mif_type_reg_w_lg_w_q_range492w493w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_mif_type_reg_w575w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_mif_type_reg_w_lg_w_lg_w_lg_w_q_range492w571w572w573w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_mif_type_reg_w_lg_w_lg_w_q_range492w571w572w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_mif_type_reg_w_lg_w_q_range492w571w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_mif_type_reg_w_q_range504w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_mif_type_reg_w_q_range499w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_mif_type_reg_w_q_range495w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_mif_type_reg_w_q_range492w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 reconf_mode_sel_reg	:	STD_LOGIC_VECTOR(2 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF reconf_mode_sel_reg : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL	 wire_reconf_mode_sel_reg_ena	:	STD_LOGIC_VECTOR(2 DOWNTO 0);
	 SIGNAL	 reconfig_data_reg	:	STD_LOGIC_VECTOR(15 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF reconfig_data_reg : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL	 wire_reconfig_data_reg_ena	:	STD_LOGIC_VECTOR(15 DOWNTO 0);
	 SIGNAL  wire_reconfig_data_reg_w_lg_w_lg_w_q_range259w476w477w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_reconfig_data_reg_w_lg_w_q_range259w476w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_reconfig_data_reg_w_lg_w_lg_w_lg_w_q_range259w476w477w478w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_reconfig_data_reg_w_q_range323w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_reconfig_data_reg_w_q_range228w	:	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  wire_reconfig_data_reg_w_q_range308w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_reconfig_data_reg_w_q_range253w	:	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  wire_reconfig_data_reg_w_q_range220w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_reconfig_data_reg_w_q_range236w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_reconfig_data_reg_w_q_range204w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_reconfig_data_reg_w_q_range259w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_reconfig_data_reg_w_q_range211w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_reconfig_data_reg_w_q_range269w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_reconfig_data_reg_w_q_range244w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_reconfig_data_reg_w_q_range314w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_reconfig_data_reg_w_q_range278w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_reconfig_data_reg_w_q_range299w	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL	 reconfig_done_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF reconfig_done_reg : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL	 wire_reconfig_done_reg_ena	:	STD_LOGIC;
	 SIGNAL  wire_reconfig_done_reg_w_lg_q468w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_reconfig_done_reg_w_lg_q469w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 state_mc_reg	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF state_mc_reg : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL	 wr_addr_inc_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF wr_addr_inc_reg : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL	 wr_rd_pulse_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF wr_rd_pulse_reg : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL	 wire_wr_rd_pulse_reg_ena	:	STD_LOGIC;
	 SIGNAL	 wire_wr_rd_pulse_reg_sclr	:	STD_LOGIC;
	 SIGNAL  wire_wr_rd_pulse_reg_w_lg_q179w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_wr_rd_pulse_reg_w_lg_q128w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 wren_data_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF wren_data_reg : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL	 wire_wren_data_reg_clrn	:	STD_LOGIC;
	 SIGNAL	 wire_wren_data_reg_ena	:	STD_LOGIC;
	 SIGNAL  wire_wren_data_reg_w_lg_q608w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_add_sub6_w_lg_w_lg_result531w532w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_add_sub6_w_lg_result531w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_add_sub6_result	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_dprio_addr_offset_cmpr_aeb	:	STD_LOGIC;
	 SIGNAL  wire_dprio_addr_offset_cmpr_datab	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_is_central_pcs490w543w544w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_is_rcxpat_chnl_en_ch_word_aeb	:	STD_LOGIC;
	 SIGNAL  wire_is_rcxpat_chnl_en_ch_word_datab	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_is_second_mif_header_address_aeb	:	STD_LOGIC;
	 SIGNAL  wire_is_second_mif_header_address_datab	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_is_special_address_aeb	:	STD_LOGIC;
	 SIGNAL  wire_is_special_address_datab	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_is_table_33_idx_aeb	:	STD_LOGIC;
	 SIGNAL  wire_is_table_33_idx_datab	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_is_table_34_idx_aeb	:	STD_LOGIC;
	 SIGNAL  wire_is_table_34_idx_datab	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_is_table_35_cmp_aeb	:	STD_LOGIC;
	 SIGNAL  wire_is_table_35_cmp_datab	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_is_table_37_cmp_aeb	:	STD_LOGIC;
	 SIGNAL  wire_is_table_37_cmp_datab	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_is_table_38_cmp_aeb	:	STD_LOGIC;
	 SIGNAL  wire_is_table_38_cmp_datab	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_is_table_42_cmp_aeb	:	STD_LOGIC;
	 SIGNAL  wire_is_table_42_cmp_datab	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_is_table_43_cmp_aeb	:	STD_LOGIC;
	 SIGNAL  wire_is_table_43_cmp_datab	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_is_table_44_cmp_aeb	:	STD_LOGIC;
	 SIGNAL  wire_is_table_44_cmp_datab	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_is_table_46_cmp_aeb	:	STD_LOGIC;
	 SIGNAL  wire_is_table_46_cmp_datab	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_is_table_47_cmp_aeb	:	STD_LOGIC;
	 SIGNAL  wire_is_table_47_cmp_datab	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_is_table_75_idx_aeb	:	STD_LOGIC;
	 SIGNAL  wire_is_table_75_idx_datab	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_is_table_76_idx_aeb	:	STD_LOGIC;
	 SIGNAL  wire_is_table_76_idx_datab	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_is_table_77_idx_aeb	:	STD_LOGIC;
	 SIGNAL  wire_is_table_77_idx_datab	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_is_table_8_idx_ageb	:	STD_LOGIC;
	 SIGNAL  wire_is_table_8_idx_datab	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_max_oper_limit_aeb	:	STD_LOGIC;
	 SIGNAL  wire_dprio_addr_offset_cnt_data	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_dprio_addr_offset_cnt_q	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_dprio_addr_offset_cnt_sclr	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_clr_offset511w512w513w514w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_mif_addr_cntr_w_lg_w_lg_q416w417w	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_mif_addr_cntr_w_lg_q416w	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_mif_addr_cntr_cnt_en	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_w_lg_en_mif_addr_cntr397w398w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_mif_addr_cntr_data	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_mif_addr_cntr_q	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_mif_addr_cntr_sclr	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_w412w413w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_mif_addr_cntr_sload	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_w_lg_w_lg_is_second_mif_header399w400w401w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_oper_count_q	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_oper_count_sclr	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_idle_state30w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_reconf_mode_dec_enable	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_w_lg_idle_state31w199w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_reconf_mode_dec_eq	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_data	:	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_result	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_central_pcs_first_word_mux_sel	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_data	:	STD_LOGIC_VECTOR (19 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_result	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_max_word_per_mif_type_sel	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_header_proc118w160w161w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_is_rcxpat_chnl_en_ch171w172w315w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_load_mif_header479w480w484w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_load_mif_header479w480w488w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_load_mif_header479w480w481w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_load_mif_header479w480w486w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_dprio_datain611w612w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_dprio_pulse600w628w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_central_pcs569w570w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_mif_header465w466w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_rcxpat_chnl_en_ch316w317w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_rx_mif_type661w662w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_tier_1175w177w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_write_reconfig_addr119w120w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_write_state384w385w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_write_word_done633w634w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_is_mif_header190w191w192w193w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_is_rx_pma515w516w518w519w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_cal_busy39w52w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_cal_busy39w45w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_cal_busy39w40w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_cal_busy39w58w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_header_proc118w160w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_analog_control113w114w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_central_pcs490w543w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_rcxpat_chnl_en_ch171w172w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_mif_header479w480w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_mif_reconfig_done389w415w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_mif_rx_only562w563w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_tx_reconfig21w22w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_write_skip170w324w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_write_skip170w229w	:	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_write_skip170w309w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_write_skip170w254w	:	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_write_skip170w221w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_write_skip170w237w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_write_skip170w290w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_write_skip170w260w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_write_skip170w212w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_write_skip170w270w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_write_skip170w245w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_write_skip170w279w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_write_skip170w300w	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w25w26w27w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_read_address115w116w117w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_write_address121w122w123w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w25w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w621w622w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_is_rx_pma515w516w517w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_is_rx_pma525w526w527w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_mif_header190w191w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_tier_1613w614w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_cal_busy41w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_w_lg_cal_busy60w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_cal_busy54w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_cal_busy47w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_clr_offset474w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_w_lg_delay_second_mif_head_out144w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_dprio_datain611w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_dprio_datain_64_67616w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_dprio_datain_68_6B615w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_dprio_datain_preemp1t617w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_dprio_datain_vodctrl618w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_dprio_pulse139w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_dprio_pulse600w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_idle_state200w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_idle_state327w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_analog_control17w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_central_pcs402w	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_central_pcs542w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_central_pcs524w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_central_pcs569w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_channel_reconfig491w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_illegal_reg_d35w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_mif_header465w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_pma_mif_type664w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_rcxpat_chnl_en_ch316w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_rx_mif_type661w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_table_33369w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_table_34529w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_table_35368w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_table_37364w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_table_38363w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_table_42362w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_table_43361w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_table_44360w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_table_46359w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_table_47358w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_table_75367w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_table_76366w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_table_77365w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_tier_1175w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_tier_1136w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_tier_1157w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_merged_dprioin357w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_mif_rx_only561w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_address115w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_wr_pulse609w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_address121w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_reconfig_addr119w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_skip322w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_skip227w	:	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_skip307w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_skip252w	:	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_skip219w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_skip235w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_skip289w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_skip258w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_skip210w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_skip268w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_skip243w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_skip313w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_skip277w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_skip298w	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_state162w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_state181w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_state448w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_state457w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_state384w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_word_done633w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_channel_address_out_range666w667w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_is_mif_header190w191w192w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w355w356w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_is_rx_pma515w516w518w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_bonded_skip169w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_cal_busy39w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_clr_offset475w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_dprio_pulse146w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_header_proc118w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_idle_state31w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_analog_control113w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_central_pcs490w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_end_mif414w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_illegal_reg_d163w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_illegal_reg_out34w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_mif_stage461w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_protected_bit168w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_rcxpat_chnl_en_ch171w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_rx_pcs498w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_table_34530w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_tier_1137w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_tx_pcs494w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_tx_pma503w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_mif_header479w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_mif_reconfig_done389w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_mif_rx_only562w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_rd_pulse73w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_state130w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_reconf_done_reg_out388w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_reset_reconf_addr159w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_reset_system447w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_rx_reconfig20w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_s0_to_08w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_s0_to_19w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_s2_to_010w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_tx_reconfig21w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_wr_pulse74w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_done19w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_mif_word_done201w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_skip170w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_state464w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_is_mif_header465w466w467w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_is_rcxpat_chnl_en_ch316w317w318w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_mif_rx_only562w563w564w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_tx_reconfig21w22w23w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_write_skip170w324w325w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_write_skip170w229w230w	:	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_write_skip170w309w310w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_write_skip170w254w255w	:	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_write_skip170w221w222w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_write_skip170w237w238w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_write_skip170w290w291w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_write_skip170w260w261w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_write_skip170w212w213w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_write_skip170w270w271w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_write_skip170w245w246w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_write_skip170w279w280w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_write_skip170w300w301w	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_w_lg_w25w26w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_cal_busy41w42w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_cal_busy60w61w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_cal_busy54w55w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_cal_busy47w48w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_dprio_datain_vodctrl618w619w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_address115w116w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_write_address121w122w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_tier_1137w178w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_tier_1137w138w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_tier_1137w158w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w319w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_tx_reconfig21w22w23w24w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_dprio_datain_vodctrl618w619w620w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w621w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w355w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w_lg_w349w350w351w352w353w354w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w349w350w351w352w353w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w349w350w351w352w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w349w350w351w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w349w350w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w134w135w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w349w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w134w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_is_table_33333w346w347w348w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_is_rcxpat_chnl_en_ch131w155w156w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_is_rcxpat_chnl_en_ch131w132w133w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_is_table_33333w346w347w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_write_skip141w142w143w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_delay_mif_head_out630w631w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_rcxpat_chnl_en_ch131w155w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_rcxpat_chnl_en_ch131w132w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_rx_pma515w516w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_rx_pma525w526w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_table_33333w346w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_write_skip141w142w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_delay_mif_head_out145w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_delay_mif_head_out630w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_mif_header190w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_rcxpat_chnl_en_ch131w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_rx_pma515w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_rx_pma525w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_table_33333w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_table_35648w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_tier_1613w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_tier_218w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_mif_header473w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_skip141w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_channel_address_range50w51w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_channel_address_out_range669w670w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  a2gr_dprio_addr :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  a2gr_dprio_data :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  a2gr_dprio_rden :	STD_LOGIC;
	 SIGNAL  a2gr_dprio_wren :	STD_LOGIC;
	 SIGNAL  a2gr_dprio_wren_data :	STD_LOGIC;
	 SIGNAL  add_sub_datab :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  add_sub_sel :	STD_LOGIC;
	 SIGNAL  bonded_skip :	STD_LOGIC;
	 SIGNAL  busy_state :	STD_LOGIC;
	 SIGNAL  cal_busy :	STD_LOGIC;
	 SIGNAL  cal_channel_address :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  cal_channel_address_out :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  cal_dprio_address :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  cal_dprioout_wire :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  cal_quad_address :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  cal_testbuses :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  central_pcs_first_word_addr :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  central_pcs_max :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  central_pcs_minus_one :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  channel_address :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  channel_address_out :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  clr_offset :	STD_LOGIC;
	 SIGNAL  default_max_limit_wire :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  delay_mif_head_out :	STD_LOGIC;
	 SIGNAL  delay_second_mif_head_out :	STD_LOGIC;
	 SIGNAL  dprio_addr_index :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  dprio_addr_offset_cnt_out :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  dprio_addr_translated_offset :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  dprio_datain :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  dprio_datain_64_67 :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  dprio_datain_68_6B :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  dprio_datain_preemp1t :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  dprio_datain_vodctrl :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  dprio_pulse :	STD_LOGIC;
	 SIGNAL  dprio_wr_done :	STD_LOGIC;
	 SIGNAL  en_mif_addr_cntr :	STD_LOGIC;
	 SIGNAL  en_write_trigger :	STD_LOGIC
	 -- synopsys translate_off
	  := '1'
	 -- synopsys translate_on
	 ;
	 SIGNAL  header_proc :	STD_LOGIC;
	 SIGNAL  idle_state :	STD_LOGIC;
	 SIGNAL  invalid_eq_dcgain :	STD_LOGIC;
	 SIGNAL  is_ageb_table_7 :	STD_LOGIC;
	 SIGNAL  is_analog_control :	STD_LOGIC;
	 SIGNAL  is_bonded_reconfig :	STD_LOGIC;
	 SIGNAL  is_cent_clk_div :	STD_LOGIC;
	 SIGNAL  is_central_pcs :	STD_LOGIC;
	 SIGNAL  is_channel_reconfig :	STD_LOGIC;
	 SIGNAL  is_end_mif :	STD_LOGIC;
	 SIGNAL  is_illegal_reg_d :	STD_LOGIC;
	 SIGNAL  is_illegal_reg_out :	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  is_mif_header :	STD_LOGIC;
	 SIGNAL  is_mif_stage :	STD_LOGIC;
	 SIGNAL  is_offset_end :	STD_LOGIC;
	 SIGNAL  is_pma_mif_type :	STD_LOGIC;
	 SIGNAL  is_protected_bit :	STD_LOGIC;
	 SIGNAL  is_rcxpat_chnl_en_ch :	STD_LOGIC;
	 SIGNAL  is_rx_mif_type :	STD_LOGIC;
	 SIGNAL  is_rx_pcs :	STD_LOGIC;
	 SIGNAL  is_rx_pma :	STD_LOGIC;
	 SIGNAL  is_second_mif_header :	STD_LOGIC;
	 SIGNAL  is_table_33 :	STD_LOGIC;
	 SIGNAL  is_table_34 :	STD_LOGIC;
	 SIGNAL  is_table_35 :	STD_LOGIC;
	 SIGNAL  is_table_37 :	STD_LOGIC;
	 SIGNAL  is_table_38 :	STD_LOGIC;
	 SIGNAL  is_table_42 :	STD_LOGIC;
	 SIGNAL  is_table_43 :	STD_LOGIC;
	 SIGNAL  is_table_44 :	STD_LOGIC;
	 SIGNAL  is_table_46 :	STD_LOGIC;
	 SIGNAL  is_table_47 :	STD_LOGIC;
	 SIGNAL  is_table_59 :	STD_LOGIC;
	 SIGNAL  is_table_61 :	STD_LOGIC;
	 SIGNAL  is_table_75 :	STD_LOGIC;
	 SIGNAL  is_table_76 :	STD_LOGIC;
	 SIGNAL  is_table_77 :	STD_LOGIC;
	 SIGNAL  is_tier_1 :	STD_LOGIC;
	 SIGNAL  is_tier_2 :	STD_LOGIC;
	 SIGNAL  is_tx_pcs :	STD_LOGIC;
	 SIGNAL  is_tx_pma :	STD_LOGIC;
	 SIGNAL  load_mif_header :	STD_LOGIC;
	 SIGNAL  merged_dprioin :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  mif_family_error :	STD_LOGIC;
	 SIGNAL  mif_reconfig_done :	STD_LOGIC;
	 SIGNAL  mif_rx_only :	STD_LOGIC;
	 SIGNAL  mif_type_error :	STD_LOGIC;
	 SIGNAL  offset_cancellation_reset	:	STD_LOGIC;
	 SIGNAL  quad_address :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  quad_address_out :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  rd_pulse :	STD_LOGIC;
	 SIGNAL  read_address :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  read_reconfig_addr :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  read_state :	STD_LOGIC;
	 SIGNAL  reconf_done_reg_out :	STD_LOGIC;
	 SIGNAL  reconfig_datain :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  reconfig_reset_all :	STD_LOGIC;
	 SIGNAL  reset_addr_done :	STD_LOGIC;
	 SIGNAL  reset_reconf_addr :	STD_LOGIC;
	 SIGNAL  reset_system :	STD_LOGIC;
	 SIGNAL  rx_pcs_max :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  rx_pma_max :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  rx_pma_minus_one :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  rx_reconfig :	STD_LOGIC;
	 SIGNAL  s0_to_0 :	STD_LOGIC;
	 SIGNAL  s0_to_1 :	STD_LOGIC;
	 SIGNAL  s0_to_2 :	STD_LOGIC;
	 SIGNAL  s2_to_0 :	STD_LOGIC;
	 SIGNAL  state_mc_reg_in :	STD_LOGIC_VECTOR (0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  table_33_data :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  table_34_addr :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  table_35_data :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  table_37_data :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  table_38_data :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  table_42_data :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  table_43_data :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  table_44_data :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  table_46_data :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  table_47_data :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  table_75_data :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  table_76_data :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  table_77_data :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  tx_pcs_max :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  tx_pma_max :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  tx_reconfig :	STD_LOGIC;
	 SIGNAL  wr_pulse :	STD_LOGIC;
	 SIGNAL  write_address :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  write_all_int :	STD_LOGIC;
	 SIGNAL  write_done :	STD_LOGIC;
	 SIGNAL  write_happened :	STD_LOGIC;
	 SIGNAL  write_mif_word_done :	STD_LOGIC;
	 SIGNAL  write_reconfig_addr :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  write_skip :	STD_LOGIC;
	 SIGNAL  write_state :	STD_LOGIC;
	 SIGNAL  write_word_64_67_data_valid :	STD_LOGIC;
	 SIGNAL  write_word_68_6B_data_valid :	STD_LOGIC;
	 SIGNAL  write_word_done :	STD_LOGIC;
	 SIGNAL  write_word_preemp1t_data_valid :	STD_LOGIC;
	 SIGNAL  write_word_vodctrl_data_valid :	STD_LOGIC;
	 SIGNAL  wire_w_cal_channel_address_range59w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_cal_channel_address_range53w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_cal_channel_address_range46w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_channel_address_range57w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_channel_address_range50w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_channel_address_out_range666w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_channel_address_out_range669w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dprio_addr_index_range647w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 COMPONENT  alt_cal_c3gxb
	 GENERIC 
	 (
		CHANNEL_ADDRESS_WIDTH	:	NATURAL := 1;
		NUMBER_OF_CHANNELS	:	NATURAL;
		SIM_MODEL_MODE	:	STRING := "FALSE";
		lpm_type	:	STRING := "alt_cal_c3gxb"
	 );
	 PORT
	 ( 
		busy	:	OUT STD_LOGIC;
		cal_error	:	OUT STD_LOGIC_VECTOR(NUMBER_OF_CHANNELS-1 DOWNTO 0);
		clock	:	IN STD_LOGIC;
		dprio_addr	:	OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		dprio_busy	:	IN STD_LOGIC;
		dprio_datain	:	IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		dprio_dataout	:	OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		dprio_rden	:	OUT STD_LOGIC;
		dprio_wren	:	OUT STD_LOGIC;
		quad_addr	:	OUT STD_LOGIC_VECTOR(8 DOWNTO 0);
		remap_addr	:	IN STD_LOGIC_VECTOR(11 DOWNTO 0) := (OTHERS => '0');
		reset	:	IN STD_LOGIC := '0';
		retain_addr	:	OUT STD_LOGIC;
		start	:	IN STD_LOGIC := '0';
		testbuses	:	IN STD_LOGIC_VECTOR(NUMBER_OF_CHANNELS-1 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
	 COMPONENT  ALTGX_RECONFIG_CIV_alt_dprio_q9l
	 PORT
	 ( 
		address	:	IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
		busy	:	OUT  STD_LOGIC;
		datain	:	IN  STD_LOGIC_VECTOR(15 DOWNTO 0) := (OTHERS => '0');
		dataout	:	OUT  STD_LOGIC_VECTOR(15 DOWNTO 0);
		dpclk	:	IN  STD_LOGIC;
		dpriodisable	:	OUT  STD_LOGIC;
		dprioin	:	OUT  STD_LOGIC;
		dprioload	:	OUT  STD_LOGIC;
		dprioout	:	IN  STD_LOGIC;
		quad_address	:	IN  STD_LOGIC_VECTOR(8 DOWNTO 0);
		rden	:	IN  STD_LOGIC := '0';
		reset	:	IN  STD_LOGIC := '0';
		status_out	:	OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		wren	:	IN  STD_LOGIC := '0';
		wren_data	:	IN  STD_LOGIC := '0'
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_add_sub
	 GENERIC 
	 (
		LPM_DIRECTION	:	STRING := "DEFAULT";
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "SIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_add_sub"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		add_sub	:	IN STD_LOGIC := '1';
		cin	:	IN STD_LOGIC := 'Z';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		cout	:	OUT STD_LOGIC;
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_compare
	 GENERIC 
	 (
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "UNSIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_compare"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		aeb	:	OUT STD_LOGIC;
		agb	:	OUT STD_LOGIC;
		ageb	:	OUT STD_LOGIC;
		alb	:	OUT STD_LOGIC;
		aleb	:	OUT STD_LOGIC;
		aneb	:	OUT STD_LOGIC;
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_counter
	 GENERIC 
	 (
		lpm_avalue	:	STRING := "0";
		lpm_direction	:	STRING := "DEFAULT";
		lpm_modulus	:	NATURAL := 0;
		lpm_port_updown	:	STRING := "PORT_CONNECTIVITY";
		lpm_pvalue	:	STRING := "0";
		lpm_svalue	:	STRING := "0";
		lpm_width	:	NATURAL;
		lpm_type	:	STRING := "lpm_counter"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		aload	:	IN STD_LOGIC := '0';
		aset	:	IN STD_LOGIC := '0';
		cin	:	IN STD_LOGIC := '1';
		clk_en	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC;
		cnt_en	:	IN STD_LOGIC := '1';
		cout	:	OUT STD_LOGIC;
		data	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		eq	:	OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		q	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0);
		sclr	:	IN STD_LOGIC := '0';
		sload	:	IN STD_LOGIC := '0';
		sset	:	IN STD_LOGIC := '0';
		updown	:	IN STD_LOGIC := '1'
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_decode
	 GENERIC 
	 (
		LPM_DECODES	:	NATURAL;
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_decode"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		data	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		enable	:	IN STD_LOGIC := '1';
		eq	:	OUT STD_LOGIC_VECTOR(LPM_DECODES-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  ALTGX_RECONFIG_CIV_mux_cda
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(35 DOWNTO 0) := (OTHERS => '0');
		result	:	OUT  STD_LOGIC_VECTOR(5 DOWNTO 0);
		sel	:	IN  STD_LOGIC_VECTOR(2 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
	 COMPONENT  ALTGX_RECONFIG_CIV_mux_8da
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(19 DOWNTO 0) := (OTHERS => '0');
		result	:	OUT  STD_LOGIC_VECTOR(4 DOWNTO 0);
		sel	:	IN  STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
 BEGIN

	wire_w_lg_w_lg_w_lg_header_proc118w160w161w(0) <= wire_w_lg_w_lg_header_proc118w160w(0) AND wire_w_lg_w_lg_is_tier_1137w158w(0);
	loop1 : FOR i IN 0 TO 1 GENERATE 
		wire_w_lg_w_lg_w_lg_is_rcxpat_chnl_en_ch171w172w315w(i) <= wire_w_lg_w_lg_is_rcxpat_chnl_en_ch171w172w(0) AND wire_reconfig_data_reg_w_q_range314w(i);
	END GENERATE loop1;
	wire_w_lg_w_lg_w_lg_load_mif_header479w480w484w(0) <= wire_w_lg_w_lg_load_mif_header479w480w(0) AND is_rx_pcs;
	wire_w_lg_w_lg_w_lg_load_mif_header479w480w488w(0) <= wire_w_lg_w_lg_load_mif_header479w480w(0) AND is_rx_pma;
	wire_w_lg_w_lg_w_lg_load_mif_header479w480w481w(0) <= wire_w_lg_w_lg_load_mif_header479w480w(0) AND is_tx_pcs;
	wire_w_lg_w_lg_w_lg_load_mif_header479w480w486w(0) <= wire_w_lg_w_lg_load_mif_header479w480w(0) AND is_tx_pma;
	loop2 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_w_lg_dprio_datain611w612w(i) <= wire_w_lg_dprio_datain611w(i) AND write_state;
	END GENERATE loop2;
	wire_w_lg_w_lg_dprio_pulse600w628w(0) <= wire_w_lg_dprio_pulse600w(0) AND is_tier_2;
	wire_w_lg_w_lg_is_central_pcs569w570w(0) <= wire_w_lg_is_central_pcs569w(0) AND dprio_pulse;
	wire_w_lg_w_lg_is_mif_header465w466w(0) <= wire_w_lg_is_mif_header465w(0) AND is_tier_1;
	loop3 : FOR i IN 0 TO 1 GENERATE 
		wire_w_lg_w_lg_is_rcxpat_chnl_en_ch316w317w(i) <= wire_w_lg_is_rcxpat_chnl_en_ch316w(0) AND wire_dprio_dataout_reg_w_q_range312w(i);
	END GENERATE loop3;
	wire_w_lg_w_lg_is_rx_mif_type661w662w(0) <= wire_w_lg_is_rx_mif_type661w(0) AND wire_w_lg_is_table_34530w(0);
	wire_w_lg_w_lg_is_tier_1175w177w(0) <= wire_w_lg_is_tier_1175w(0) AND wire_w_lg_w_lg_w_lg_is_rcxpat_chnl_en_ch131w155w156w(0);
	loop4 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_w_lg_write_reconfig_addr119w120w(i) <= wire_w_lg_write_reconfig_addr119w(i) AND wire_w_lg_header_proc118w(0);
	END GENERATE loop4;
	wire_w_lg_w_lg_write_state384w385w(0) <= wire_w_lg_write_state384w(0) AND write_happened;
	wire_w_lg_w_lg_write_word_done633w634w(0) <= wire_w_lg_write_word_done633w(0) AND is_analog_control;
	wire_w_lg_w_lg_w_lg_w_lg_is_mif_header190w191w192w193w(0) <= wire_w_lg_w_lg_w_lg_is_mif_header190w191w192w(0) AND mif_stage;
	loop5 : FOR i IN 0 TO 4 GENERATE 
		wire_w_lg_w_lg_w_lg_w_lg_is_rx_pma515w516w518w519w(i) <= wire_w_lg_w_lg_w_lg_is_rx_pma515w516w518w(0) AND wire_dprio_addr_offset_cnt_q(i);
	END GENERATE loop5;
	wire_w_lg_w_lg_cal_busy39w52w(0) <= wire_w_lg_cal_busy39w(0) AND wire_w_lg_w_channel_address_range50w51w(0);
	wire_w_lg_w_lg_cal_busy39w45w(0) <= wire_w_lg_cal_busy39w(0) AND is_central_pcs;
	loop6 : FOR i IN 0 TO 8 GENERATE 
		wire_w_lg_w_lg_cal_busy39w40w(i) <= wire_w_lg_cal_busy39w(0) AND quad_address(i);
	END GENERATE loop6;
	wire_w_lg_w_lg_cal_busy39w58w(0) <= wire_w_lg_cal_busy39w(0) AND wire_w_channel_address_range57w(0);
	wire_w_lg_w_lg_header_proc118w160w(0) <= wire_w_lg_header_proc118w(0) AND wire_w_lg_reset_reconf_addr159w(0);
	loop7 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_w_lg_is_analog_control113w114w(i) <= wire_w_lg_is_analog_control113w(0) AND read_reconfig_addr(i);
	END GENERATE loop7;
	loop8 : FOR i IN 0 TO 4 GENERATE 
		wire_w_lg_w_lg_is_central_pcs490w543w(i) <= wire_w_lg_is_central_pcs490w(0) AND wire_max_word_per_mif_type_result(i);
	END GENERATE loop8;
	wire_w_lg_w_lg_is_rcxpat_chnl_en_ch171w172w(0) <= wire_w_lg_is_rcxpat_chnl_en_ch171w(0) AND wire_w_lg_write_skip170w(0);
	wire_w_lg_w_lg_load_mif_header479w480w(0) <= wire_w_lg_load_mif_header479w(0) AND clr_offset;
	wire_w_lg_w_lg_mif_reconfig_done389w415w(0) <= wire_w_lg_mif_reconfig_done389w(0) AND wire_w_lg_is_end_mif414w(0);
	wire_w_lg_w_lg_mif_rx_only562w563w(0) <= wire_w_lg_mif_rx_only562w(0) AND wire_mif_type_reg_w_q_range499w(0);
	wire_w_lg_w_lg_tx_reconfig21w22w(0) <= wire_w_lg_tx_reconfig21w(0) AND wire_w_lg_rx_reconfig20w(0);
	wire_w_lg_w_lg_write_skip170w324w(0) <= wire_w_lg_write_skip170w(0) AND wire_reconfig_data_reg_w_q_range323w(0);
	loop9 : FOR i IN 0 TO 10 GENERATE 
		wire_w_lg_w_lg_write_skip170w229w(i) <= wire_w_lg_write_skip170w(0) AND wire_reconfig_data_reg_w_q_range228w(i);
	END GENERATE loop9;
	loop10 : FOR i IN 0 TO 8 GENERATE 
		wire_w_lg_w_lg_write_skip170w309w(i) <= wire_w_lg_write_skip170w(0) AND wire_reconfig_data_reg_w_q_range308w(i);
	END GENERATE loop10;
	loop11 : FOR i IN 0 TO 13 GENERATE 
		wire_w_lg_w_lg_write_skip170w254w(i) <= wire_w_lg_write_skip170w(0) AND wire_reconfig_data_reg_w_q_range253w(i);
	END GENERATE loop11;
	loop12 : FOR i IN 0 TO 1 GENERATE 
		wire_w_lg_w_lg_write_skip170w221w(i) <= wire_w_lg_write_skip170w(0) AND wire_reconfig_data_reg_w_q_range220w(i);
	END GENERATE loop12;
	loop13 : FOR i IN 0 TO 8 GENERATE 
		wire_w_lg_w_lg_write_skip170w237w(i) <= wire_w_lg_write_skip170w(0) AND wire_reconfig_data_reg_w_q_range236w(i);
	END GENERATE loop13;
	loop14 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_w_lg_write_skip170w290w(i) <= wire_w_lg_write_skip170w(0) AND wire_reconfig_data_reg_w_q_range204w(i);
	END GENERATE loop14;
	loop15 : FOR i IN 0 TO 3 GENERATE 
		wire_w_lg_w_lg_write_skip170w260w(i) <= wire_w_lg_write_skip170w(0) AND wire_reconfig_data_reg_w_q_range259w(i);
	END GENERATE loop15;
	wire_w_lg_w_lg_write_skip170w212w(0) <= wire_w_lg_write_skip170w(0) AND wire_reconfig_data_reg_w_q_range211w(0);
	loop16 : FOR i IN 0 TO 8 GENERATE 
		wire_w_lg_w_lg_write_skip170w270w(i) <= wire_w_lg_write_skip170w(0) AND wire_reconfig_data_reg_w_q_range269w(i);
	END GENERATE loop16;
	loop17 : FOR i IN 0 TO 2 GENERATE 
		wire_w_lg_w_lg_write_skip170w245w(i) <= wire_w_lg_write_skip170w(0) AND wire_reconfig_data_reg_w_q_range244w(i);
	END GENERATE loop17;
	loop18 : FOR i IN 0 TO 4 GENERATE 
		wire_w_lg_w_lg_write_skip170w279w(i) <= wire_w_lg_write_skip170w(0) AND wire_reconfig_data_reg_w_q_range278w(i);
	END GENERATE loop18;
	loop19 : FOR i IN 0 TO 9 GENERATE 
		wire_w_lg_w_lg_write_skip170w300w(i) <= wire_w_lg_write_skip170w(0) AND wire_reconfig_data_reg_w_q_range299w(i);
	END GENERATE loop19;
	wire_w_lg_w_lg_w25w26w27w(0) <= wire_w_lg_w25w26w(0) AND write_state;
	loop20 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_w_lg_w_lg_read_address115w116w117w(i) <= wire_w_lg_w_lg_read_address115w116w(i) AND read_state;
	END GENERATE loop20;
	loop21 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_w_lg_w_lg_write_address121w122w123w(i) <= wire_w_lg_w_lg_write_address121w122w(i) AND write_state;
	END GENERATE loop21;
	wire_w25w(0) <= wire_w_lg_w_lg_w_lg_w_lg_tx_reconfig21w22w23w24w(0) AND is_tier_1;
	loop22 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_w621w622w(i) <= wire_w621w(i) AND is_analog_control;
	END GENERATE loop22;
	loop23 : FOR i IN 0 TO 4 GENERATE 
		wire_w_lg_w_lg_w_lg_is_rx_pma515w516w517w(i) <= wire_w_lg_w_lg_is_rx_pma515w516w(0) AND dprio_addr_translated_offset(i);
	END GENERATE loop23;
	loop24 : FOR i IN 0 TO 4 GENERATE 
		wire_w_lg_w_lg_w_lg_is_rx_pma525w526w527w(i) <= wire_w_lg_w_lg_is_rx_pma525w526w(0) AND rx_pma_minus_one(i);
	END GENERATE loop24;
	wire_w_lg_w_lg_is_mif_header190w191w(0) <= wire_w_lg_is_mif_header190w(0) AND dprio_pulse;
	loop25 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_w_lg_is_tier_1613w614w(i) <= wire_w_lg_is_tier_1613w(0) AND reconfig_datain(i);
	END GENERATE loop25;
	loop26 : FOR i IN 0 TO 8 GENERATE 
		wire_w_lg_cal_busy41w(i) <= cal_busy AND cal_quad_address(i);
	END GENERATE loop26;
	wire_w_lg_cal_busy60w(0) <= cal_busy AND wire_w_cal_channel_address_range59w(0);
	wire_w_lg_cal_busy54w(0) <= cal_busy AND wire_w_cal_channel_address_range53w(0);
	wire_w_lg_cal_busy47w(0) <= cal_busy AND wire_w_cal_channel_address_range46w(0);
	loop27 : FOR i IN 0 TO 3 GENERATE 
		wire_w_lg_clr_offset474w(i) <= clr_offset AND mif_type_reg(i);
	END GENERATE loop27;
	wire_w_lg_delay_second_mif_head_out144w(0) <= delay_second_mif_head_out AND wire_w_lg_w_lg_w_lg_write_skip141w142w143w(0);
	loop28 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_dprio_datain611w(i) <= dprio_datain(i) AND wire_w_lg_header_proc118w(0);
	END GENERATE loop28;
	loop29 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_dprio_datain_64_67616w(i) <= dprio_datain_64_67(i) AND write_word_64_67_data_valid;
	END GENERATE loop29;
	loop30 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_dprio_datain_68_6B615w(i) <= dprio_datain_68_6B(i) AND write_word_68_6B_data_valid;
	END GENERATE loop30;
	loop31 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_dprio_datain_preemp1t617w(i) <= dprio_datain_preemp1t(i) AND write_word_preemp1t_data_valid;
	END GENERATE loop31;
	loop32 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_dprio_datain_vodctrl618w(i) <= dprio_datain_vodctrl(i) AND write_word_vodctrl_data_valid;
	END GENERATE loop32;
	wire_w_lg_dprio_pulse139w(0) <= dprio_pulse AND wire_w_lg_w_lg_is_tier_1137w138w(0);
	wire_w_lg_dprio_pulse600w(0) <= dprio_pulse AND write_happened;
	wire_w_lg_idle_state200w(0) <= idle_state AND wire_mif_stage_w_lg_q194w(0);
	wire_w_lg_idle_state327w(0) <= idle_state AND write_all;
	wire_w_lg_is_analog_control17w(0) <= is_analog_control AND write_state;
	loop33 : FOR i IN 0 TO 5 GENERATE 
		wire_w_lg_is_central_pcs402w(i) <= is_central_pcs AND central_pcs_first_word_addr(i);
	END GENERATE loop33;
	loop34 : FOR i IN 0 TO 4 GENERATE 
		wire_w_lg_is_central_pcs542w(i) <= is_central_pcs AND central_pcs_max(i);
	END GENERATE loop34;
	loop35 : FOR i IN 0 TO 4 GENERATE 
		wire_w_lg_is_central_pcs524w(i) <= is_central_pcs AND central_pcs_minus_one(i);
	END GENERATE loop35;
	wire_w_lg_is_central_pcs569w(0) <= is_central_pcs AND is_offset_end;
	wire_w_lg_is_channel_reconfig491w(0) <= is_channel_reconfig AND wire_w_lg_is_central_pcs490w(0);
	wire_w_lg_is_illegal_reg_d35w(0) <= is_illegal_reg_d AND wire_w_lg_write_done19w(0);
	wire_w_lg_is_mif_header465w(0) <= is_mif_header AND wire_w_lg_write_state464w(0);
	wire_w_lg_is_pma_mif_type664w(0) <= is_pma_mif_type AND wire_w_lg_is_central_pcs490w(0);
	wire_w_lg_is_rcxpat_chnl_en_ch316w(0) <= is_rcxpat_chnl_en_ch AND wire_w_lg_write_skip170w(0);
	wire_w_lg_is_rx_mif_type661w(0) <= is_rx_mif_type AND wire_w_lg_is_central_pcs490w(0);
	loop36 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_is_table_33369w(i) <= is_table_33 AND table_33_data(i);
	END GENERATE loop36;
	loop37 : FOR i IN 0 TO 4 GENERATE 
		wire_w_lg_is_table_34529w(i) <= is_table_34 AND table_34_addr(i);
	END GENERATE loop37;
	loop38 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_is_table_35368w(i) <= is_table_35 AND table_35_data(i);
	END GENERATE loop38;
	loop39 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_is_table_37364w(i) <= is_table_37 AND table_37_data(i);
	END GENERATE loop39;
	loop40 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_is_table_38363w(i) <= is_table_38 AND table_38_data(i);
	END GENERATE loop40;
	loop41 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_is_table_42362w(i) <= is_table_42 AND table_42_data(i);
	END GENERATE loop41;
	loop42 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_is_table_43361w(i) <= is_table_43 AND table_43_data(i);
	END GENERATE loop42;
	loop43 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_is_table_44360w(i) <= is_table_44 AND table_44_data(i);
	END GENERATE loop43;
	loop44 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_is_table_46359w(i) <= is_table_46 AND table_46_data(i);
	END GENERATE loop44;
	loop45 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_is_table_47358w(i) <= is_table_47 AND table_47_data(i);
	END GENERATE loop45;
	loop46 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_is_table_75367w(i) <= is_table_75 AND table_75_data(i);
	END GENERATE loop46;
	loop47 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_is_table_76366w(i) <= is_table_76 AND table_76_data(i);
	END GENERATE loop47;
	loop48 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_is_table_77365w(i) <= is_table_77 AND table_77_data(i);
	END GENERATE loop48;
	wire_w_lg_is_tier_1175w(0) <= is_tier_1 AND wire_w_lg_header_proc118w(0);
	wire_w_lg_is_tier_1136w(0) <= is_tier_1 AND wire_w_lg_w134w135w(0);
	wire_w_lg_is_tier_1157w(0) <= is_tier_1 AND wire_w_lg_w_lg_w_lg_is_rcxpat_chnl_en_ch131w155w156w(0);
	loop49 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_merged_dprioin357w(i) <= merged_dprioin(i) AND wire_w_lg_w355w356w(0);
	END GENERATE loop49;
	wire_w_lg_mif_rx_only561w(0) <= mif_rx_only AND wire_mif_type_reg_w_q_range492w(0);
	loop50 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_read_address115w(i) <= read_address(i) AND is_analog_control;
	END GENERATE loop50;
	wire_w_lg_wr_pulse609w(0) <= wr_pulse AND wire_wren_data_reg_w_lg_q608w(0);
	loop51 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_write_address121w(i) <= write_address(i) AND is_analog_control;
	END GENERATE loop51;
	loop52 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_write_reconfig_addr119w(i) <= write_reconfig_addr(i) AND wire_w_lg_is_analog_control113w(0);
	END GENERATE loop52;
	wire_w_lg_write_skip322w(0) <= write_skip AND wire_dprio_dataout_reg_w_q_range321w(0);
	loop53 : FOR i IN 0 TO 10 GENERATE 
		wire_w_lg_write_skip227w(i) <= write_skip AND wire_dprio_dataout_reg_w_q_range226w(i);
	END GENERATE loop53;
	loop54 : FOR i IN 0 TO 8 GENERATE 
		wire_w_lg_write_skip307w(i) <= write_skip AND wire_dprio_dataout_reg_w_q_range264w(i);
	END GENERATE loop54;
	loop55 : FOR i IN 0 TO 13 GENERATE 
		wire_w_lg_write_skip252w(i) <= write_skip AND wire_dprio_dataout_reg_w_q_range251w(i);
	END GENERATE loop55;
	loop56 : FOR i IN 0 TO 1 GENERATE 
		wire_w_lg_write_skip219w(i) <= write_skip AND wire_dprio_dataout_reg_w_q_range218w(i);
	END GENERATE loop56;
	loop57 : FOR i IN 0 TO 8 GENERATE 
		wire_w_lg_write_skip235w(i) <= write_skip AND wire_dprio_dataout_reg_w_q_range234w(i);
	END GENERATE loop57;
	loop58 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_write_skip289w(i) <= write_skip AND wire_dprio_dataout_reg_w_q_range288w(i);
	END GENERATE loop58;
	loop59 : FOR i IN 0 TO 3 GENERATE 
		wire_w_lg_write_skip258w(i) <= write_skip AND wire_dprio_dataout_reg_w_q_range257w(i);
	END GENERATE loop59;
	wire_w_lg_write_skip210w(0) <= write_skip AND wire_dprio_dataout_reg_w_q_range209w(0);
	loop60 : FOR i IN 0 TO 8 GENERATE 
		wire_w_lg_write_skip268w(i) <= write_skip AND wire_dprio_dataout_reg_w_q_range267w(i);
	END GENERATE loop60;
	loop61 : FOR i IN 0 TO 2 GENERATE 
		wire_w_lg_write_skip243w(i) <= write_skip AND wire_dprio_dataout_reg_w_q_range242w(i);
	END GENERATE loop61;
	loop62 : FOR i IN 0 TO 1 GENERATE 
		wire_w_lg_write_skip313w(i) <= write_skip AND wire_dprio_dataout_reg_w_q_range312w(i);
	END GENERATE loop62;
	loop63 : FOR i IN 0 TO 4 GENERATE 
		wire_w_lg_write_skip277w(i) <= write_skip AND wire_dprio_dataout_reg_w_q_range276w(i);
	END GENERATE loop63;
	loop64 : FOR i IN 0 TO 9 GENERATE 
		wire_w_lg_write_skip298w(i) <= write_skip AND wire_dprio_dataout_reg_w_q_range297w(i);
	END GENERATE loop64;
	wire_w_lg_write_state162w(0) <= write_state AND wire_w_lg_w_lg_w_lg_header_proc118w160w161w(0);
	wire_w_lg_write_state181w(0) <= write_state AND wire_w_lg_dprio_pulse146w(0);
	wire_w_lg_write_state448w(0) <= write_state AND wire_w_lg_reconf_done_reg_out388w(0);
	wire_w_lg_write_state457w(0) <= write_state AND wire_w_lg_write_mif_word_done201w(0);
	wire_w_lg_write_state384w(0) <= write_state AND dprio_wr_done;
	wire_w_lg_write_word_done633w(0) <= write_word_done AND write_happened;
	wire_w_lg_w_channel_address_out_range666w667w(0) <= wire_w_channel_address_out_range666w(0) AND wire_w_lg_is_central_pcs490w(0);
	wire_w_lg_w_lg_w_lg_is_mif_header190w191w192w(0) <= NOT wire_w_lg_w_lg_is_mif_header190w191w(0);
	wire_w_lg_w355w356w(0) <= NOT wire_w355w(0);
	wire_w_lg_w_lg_w_lg_is_rx_pma515w516w518w(0) <= NOT wire_w_lg_w_lg_is_rx_pma515w516w(0);
	wire_w_lg_bonded_skip169w(0) <= NOT bonded_skip;
	wire_w_lg_cal_busy39w(0) <= NOT cal_busy;
	wire_w_lg_clr_offset475w(0) <= NOT clr_offset;
	wire_w_lg_dprio_pulse146w(0) <= NOT dprio_pulse;
	wire_w_lg_header_proc118w(0) <= NOT header_proc;
	wire_w_lg_idle_state31w(0) <= NOT idle_state;
	wire_w_lg_is_analog_control113w(0) <= NOT is_analog_control;
	wire_w_lg_is_central_pcs490w(0) <= NOT is_central_pcs;
	wire_w_lg_is_end_mif414w(0) <= NOT is_end_mif;
	wire_w_lg_is_illegal_reg_d163w(0) <= NOT is_illegal_reg_d;
	wire_w_lg_is_illegal_reg_out34w(0) <= NOT is_illegal_reg_out;
	wire_w_lg_is_mif_stage461w(0) <= NOT is_mif_stage;
	wire_w_lg_is_protected_bit168w(0) <= NOT is_protected_bit;
	wire_w_lg_is_rcxpat_chnl_en_ch171w(0) <= NOT is_rcxpat_chnl_en_ch;
	wire_w_lg_is_rx_pcs498w(0) <= NOT is_rx_pcs;
	wire_w_lg_is_table_34530w(0) <= NOT is_table_34;
	wire_w_lg_is_tier_1137w(0) <= NOT is_tier_1;
	wire_w_lg_is_tx_pcs494w(0) <= NOT is_tx_pcs;
	wire_w_lg_is_tx_pma503w(0) <= NOT is_tx_pma;
	wire_w_lg_load_mif_header479w(0) <= NOT load_mif_header;
	wire_w_lg_mif_reconfig_done389w(0) <= NOT mif_reconfig_done;
	wire_w_lg_mif_rx_only562w(0) <= NOT mif_rx_only;
	wire_w_lg_rd_pulse73w(0) <= NOT rd_pulse;
	wire_w_lg_read_state130w(0) <= NOT read_state;
	wire_w_lg_reconf_done_reg_out388w(0) <= NOT reconf_done_reg_out;
	wire_w_lg_reset_reconf_addr159w(0) <= NOT reset_reconf_addr;
	wire_w_lg_reset_system447w(0) <= NOT reset_system;
	wire_w_lg_rx_reconfig20w(0) <= NOT rx_reconfig;
	wire_w_lg_s0_to_08w(0) <= NOT s0_to_0;
	wire_w_lg_s0_to_19w(0) <= NOT s0_to_1;
	wire_w_lg_s2_to_010w(0) <= NOT s2_to_0;
	wire_w_lg_tx_reconfig21w(0) <= NOT tx_reconfig;
	wire_w_lg_wr_pulse74w(0) <= NOT wr_pulse;
	wire_w_lg_write_done19w(0) <= NOT write_done;
	wire_w_lg_write_mif_word_done201w(0) <= NOT write_mif_word_done;
	wire_w_lg_write_skip170w(0) <= NOT write_skip;
	wire_w_lg_write_state464w(0) <= NOT write_state;
	wire_w_lg_w_lg_w_lg_is_mif_header465w466w467w(0) <= wire_w_lg_w_lg_is_mif_header465w466w(0) OR wire_w_lg_is_tier_1137w(0);
	loop65 : FOR i IN 0 TO 1 GENERATE 
		wire_w_lg_w_lg_w_lg_is_rcxpat_chnl_en_ch316w317w318w(i) <= wire_w_lg_w_lg_is_rcxpat_chnl_en_ch316w317w(i) OR wire_w_lg_w_lg_w_lg_is_rcxpat_chnl_en_ch171w172w315w(i);
	END GENERATE loop65;
	wire_w_lg_w_lg_w_lg_mif_rx_only562w563w564w(0) <= wire_w_lg_w_lg_mif_rx_only562w563w(0) OR wire_w_lg_mif_rx_only561w(0);
	wire_w_lg_w_lg_w_lg_tx_reconfig21w22w23w(0) <= wire_w_lg_w_lg_tx_reconfig21w22w(0) OR mif_type_error;
	wire_w_lg_w_lg_w_lg_write_skip170w324w325w(0) <= wire_w_lg_w_lg_write_skip170w324w(0) OR wire_w_lg_write_skip322w(0);
	loop66 : FOR i IN 0 TO 10 GENERATE 
		wire_w_lg_w_lg_w_lg_write_skip170w229w230w(i) <= wire_w_lg_w_lg_write_skip170w229w(i) OR wire_w_lg_write_skip227w(i);
	END GENERATE loop66;
	loop67 : FOR i IN 0 TO 8 GENERATE 
		wire_w_lg_w_lg_w_lg_write_skip170w309w310w(i) <= wire_w_lg_w_lg_write_skip170w309w(i) OR wire_w_lg_write_skip307w(i);
	END GENERATE loop67;
	loop68 : FOR i IN 0 TO 13 GENERATE 
		wire_w_lg_w_lg_w_lg_write_skip170w254w255w(i) <= wire_w_lg_w_lg_write_skip170w254w(i) OR wire_w_lg_write_skip252w(i);
	END GENERATE loop68;
	loop69 : FOR i IN 0 TO 1 GENERATE 
		wire_w_lg_w_lg_w_lg_write_skip170w221w222w(i) <= wire_w_lg_w_lg_write_skip170w221w(i) OR wire_w_lg_write_skip219w(i);
	END GENERATE loop69;
	loop70 : FOR i IN 0 TO 8 GENERATE 
		wire_w_lg_w_lg_w_lg_write_skip170w237w238w(i) <= wire_w_lg_w_lg_write_skip170w237w(i) OR wire_w_lg_write_skip235w(i);
	END GENERATE loop70;
	loop71 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_w_lg_w_lg_write_skip170w290w291w(i) <= wire_w_lg_w_lg_write_skip170w290w(i) OR wire_w_lg_write_skip289w(i);
	END GENERATE loop71;
	loop72 : FOR i IN 0 TO 3 GENERATE 
		wire_w_lg_w_lg_w_lg_write_skip170w260w261w(i) <= wire_w_lg_w_lg_write_skip170w260w(i) OR wire_w_lg_write_skip258w(i);
	END GENERATE loop72;
	wire_w_lg_w_lg_w_lg_write_skip170w212w213w(0) <= wire_w_lg_w_lg_write_skip170w212w(0) OR wire_w_lg_write_skip210w(0);
	loop73 : FOR i IN 0 TO 8 GENERATE 
		wire_w_lg_w_lg_w_lg_write_skip170w270w271w(i) <= wire_w_lg_w_lg_write_skip170w270w(i) OR wire_w_lg_write_skip268w(i);
	END GENERATE loop73;
	loop74 : FOR i IN 0 TO 2 GENERATE 
		wire_w_lg_w_lg_w_lg_write_skip170w245w246w(i) <= wire_w_lg_w_lg_write_skip170w245w(i) OR wire_w_lg_write_skip243w(i);
	END GENERATE loop74;
	loop75 : FOR i IN 0 TO 4 GENERATE 
		wire_w_lg_w_lg_w_lg_write_skip170w279w280w(i) <= wire_w_lg_w_lg_write_skip170w279w(i) OR wire_w_lg_write_skip277w(i);
	END GENERATE loop75;
	loop76 : FOR i IN 0 TO 9 GENERATE 
		wire_w_lg_w_lg_w_lg_write_skip170w300w301w(i) <= wire_w_lg_w_lg_write_skip170w300w(i) OR wire_w_lg_write_skip298w(i);
	END GENERATE loop76;
	wire_w_lg_w25w26w(0) <= wire_w25w(0) OR invalid_eq_dcgain;
	loop77 : FOR i IN 0 TO 8 GENERATE 
		wire_w_lg_w_lg_cal_busy41w42w(i) <= wire_w_lg_cal_busy41w(i) OR wire_w_lg_w_lg_cal_busy39w40w(i);
	END GENERATE loop77;
	wire_w_lg_w_lg_cal_busy60w61w(0) <= wire_w_lg_cal_busy60w(0) OR wire_w_lg_w_lg_cal_busy39w58w(0);
	wire_w_lg_w_lg_cal_busy54w55w(0) <= wire_w_lg_cal_busy54w(0) OR wire_w_lg_w_lg_cal_busy39w52w(0);
	wire_w_lg_w_lg_cal_busy47w48w(0) <= wire_w_lg_cal_busy47w(0) OR wire_w_lg_w_lg_cal_busy39w45w(0);
	loop78 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_w_lg_dprio_datain_vodctrl618w619w(i) <= wire_w_lg_dprio_datain_vodctrl618w(i) OR wire_w_lg_dprio_datain_preemp1t617w(i);
	END GENERATE loop78;
	loop79 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_w_lg_read_address115w116w(i) <= wire_w_lg_read_address115w(i) OR wire_w_lg_w_lg_is_analog_control113w114w(i);
	END GENERATE loop79;
	loop80 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_w_lg_write_address121w122w(i) <= wire_w_lg_write_address121w(i) OR wire_w_lg_w_lg_write_reconfig_addr119w120w(i);
	END GENERATE loop80;
	wire_w_lg_w_lg_is_tier_1137w178w(0) <= wire_w_lg_is_tier_1137w(0) OR wire_w_lg_w_lg_is_tier_1175w177w(0);
	wire_w_lg_w_lg_is_tier_1137w138w(0) <= wire_w_lg_is_tier_1137w(0) OR wire_w_lg_is_tier_1136w(0);
	wire_w_lg_w_lg_is_tier_1137w158w(0) <= wire_w_lg_is_tier_1137w(0) OR wire_w_lg_is_tier_1157w(0);
	loop81 : FOR i IN 0 TO 1 GENERATE 
		wire_w319w(i) <= wire_w_lg_w_lg_w_lg_is_rcxpat_chnl_en_ch316w317w318w(i) OR wire_w_lg_write_skip313w(i);
	END GENERATE loop81;
	wire_w_lg_w_lg_w_lg_w_lg_tx_reconfig21w22w23w24w(0) <= wire_w_lg_w_lg_w_lg_tx_reconfig21w22w23w(0) OR mif_family_error;
	loop82 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_w_lg_w_lg_dprio_datain_vodctrl618w619w620w(i) <= wire_w_lg_w_lg_dprio_datain_vodctrl618w619w(i) OR wire_w_lg_dprio_datain_64_67616w(i);
	END GENERATE loop82;
	loop83 : FOR i IN 0 TO 15 GENERATE 
		wire_w621w(i) <= wire_w_lg_w_lg_w_lg_dprio_datain_vodctrl618w619w620w(i) OR wire_w_lg_dprio_datain_68_6B615w(i);
	END GENERATE loop83;
	wire_w355w(0) <= wire_w_lg_w_lg_w_lg_w_lg_w_lg_w349w350w351w352w353w354w(0) OR is_table_47;
	wire_w_lg_w_lg_w_lg_w_lg_w_lg_w349w350w351w352w353w354w(0) <= wire_w_lg_w_lg_w_lg_w_lg_w349w350w351w352w353w(0) OR is_table_46;
	wire_w_lg_w_lg_w_lg_w_lg_w349w350w351w352w353w(0) <= wire_w_lg_w_lg_w_lg_w349w350w351w352w(0) OR is_table_44;
	wire_w_lg_w_lg_w_lg_w349w350w351w352w(0) <= wire_w_lg_w_lg_w349w350w351w(0) OR is_table_43;
	wire_w_lg_w_lg_w349w350w351w(0) <= wire_w_lg_w349w350w(0) OR is_table_42;
	wire_w_lg_w349w350w(0) <= wire_w349w(0) OR is_table_38;
	wire_w_lg_w134w135w(0) <= wire_w134w(0) OR is_cent_clk_div;
	wire_w349w(0) <= wire_w_lg_w_lg_w_lg_w_lg_is_table_33333w346w347w348w(0) OR is_table_37;
	wire_w134w(0) <= wire_w_lg_w_lg_w_lg_is_rcxpat_chnl_en_ch131w132w133w(0) OR is_protected_bit;
	wire_w_lg_w_lg_w_lg_w_lg_is_table_33333w346w347w348w(0) <= wire_w_lg_w_lg_w_lg_is_table_33333w346w347w(0) OR is_table_77;
	wire_w_lg_w_lg_w_lg_is_rcxpat_chnl_en_ch131w155w156w(0) <= wire_w_lg_w_lg_is_rcxpat_chnl_en_ch131w155w(0) OR is_protected_bit;
	wire_w_lg_w_lg_w_lg_is_rcxpat_chnl_en_ch131w132w133w(0) <= wire_w_lg_w_lg_is_rcxpat_chnl_en_ch131w132w(0) OR bonded_skip;
	wire_w_lg_w_lg_w_lg_is_table_33333w346w347w(0) <= wire_w_lg_w_lg_is_table_33333w346w(0) OR is_table_76;
	wire_w_lg_w_lg_w_lg_write_skip141w142w143w(0) <= wire_w_lg_w_lg_write_skip141w142w(0) OR is_cent_clk_div;
	wire_w_lg_w_lg_delay_mif_head_out630w631w(0) <= wire_w_lg_delay_mif_head_out630w(0) OR write_mif_word_done;
	wire_w_lg_w_lg_is_rcxpat_chnl_en_ch131w155w(0) <= wire_w_lg_is_rcxpat_chnl_en_ch131w(0) OR bonded_skip;
	wire_w_lg_w_lg_is_rcxpat_chnl_en_ch131w132w(0) <= wire_w_lg_is_rcxpat_chnl_en_ch131w(0) OR is_mif_header;
	wire_w_lg_w_lg_is_rx_pma515w516w(0) <= wire_w_lg_is_rx_pma515w(0) OR is_ageb_table_7;
	wire_w_lg_w_lg_is_rx_pma525w526w(0) <= wire_w_lg_is_rx_pma525w(0) OR is_ageb_table_7;
	wire_w_lg_w_lg_is_table_33333w346w(0) <= wire_w_lg_is_table_33333w(0) OR is_table_75;
	wire_w_lg_w_lg_write_skip141w142w(0) <= wire_w_lg_write_skip141w(0) OR is_protected_bit;
	wire_w_lg_delay_mif_head_out145w(0) <= delay_mif_head_out OR wire_w_lg_delay_second_mif_head_out144w(0);
	wire_w_lg_delay_mif_head_out630w(0) <= delay_mif_head_out OR delay_second_mif_head_out;
	wire_w_lg_is_mif_header190w(0) <= is_mif_header OR mif_reconfig_done;
	wire_w_lg_is_rcxpat_chnl_en_ch131w(0) <= is_rcxpat_chnl_en_ch OR write_skip;
	wire_w_lg_is_rx_pma515w(0) <= is_rx_pma OR is_central_pcs;
	wire_w_lg_is_rx_pma525w(0) <= is_rx_pma OR is_rx_pcs;
	wire_w_lg_is_table_33333w(0) <= is_table_33 OR is_table_35;
	wire_w_lg_is_table_35648w(0) <= is_table_35 OR wire_w_dprio_addr_index_range647w(0);
	wire_w_lg_is_tier_1613w(0) <= is_tier_1 OR is_tier_2;
	wire_w_lg_is_tier_218w(0) <= is_tier_2 OR wire_w_lg_is_analog_control17w(0);
	wire_w_lg_load_mif_header473w(0) <= load_mif_header OR clr_offset;
	wire_w_lg_write_skip141w(0) <= write_skip OR bonded_skip;
	wire_w_lg_w_channel_address_range50w51w(0) <= wire_w_channel_address_range50w(0) OR is_central_pcs;
	wire_w_lg_w_channel_address_out_range669w670w(0) <= wire_w_channel_address_out_range669w(0) OR is_central_pcs;
	a2gr_dprio_addr <= (wire_w_lg_w_lg_w_lg_write_address121w122w123w OR wire_w_lg_w_lg_w_lg_read_address115w116w117w);
	a2gr_dprio_data <= wire_w_lg_w_lg_dprio_datain611w612w;
	a2gr_dprio_rden <= rd_pulse;
	a2gr_dprio_wren <= (wire_w_lg_wr_pulse609w(0) AND wire_w_lg_is_analog_control113w(0));
	a2gr_dprio_wren_data <= (wr_pulse AND (wren_data_reg OR is_analog_control));
	add_sub_datab <= (wire_w_lg_w_lg_w_lg_is_rx_pma525w526w527w OR wire_w_lg_is_central_pcs524w);
	add_sub_sel <= ((NOT (wire_w_lg_is_rx_pma515w(0) OR is_rx_pcs)) OR is_ageb_table_7);
	bonded_skip <= ((((((wire_w_lg_is_table_33333w(0) AND is_bonded_reconfig) OR is_table_59) OR is_table_61) OR is_table_75) OR is_table_76) OR is_table_77);
	busy <= (busy_state OR cal_busy);
	busy_state <= (read_state OR write_state);
	cal_busy <= wire_calibration_c3gxb_busy;
	cal_channel_address <= wire_calibration_c3gxb_dprio_addr(14 DOWNTO 12);
	cal_channel_address_out <= address_pres_reg(2 DOWNTO 0);
	cal_dprio_address <= ( wire_calibration_c3gxb_dprio_addr(15) & cal_channel_address_out & wire_calibration_c3gxb_dprio_addr(11 DOWNTO 0));
	cal_dprioout_wire(0) <= ( reconfig_fromgxb(0));
	cal_quad_address <= wire_calibration_c3gxb_quad_addr;
	cal_testbuses(0) <= ( reconfig_fromgxb(1));
	central_pcs_first_word_addr <= wire_central_pcs_first_word_mux_result;
	central_pcs_max <= "00100";
	central_pcs_minus_one <= "00001";
	channel_address <= (OTHERS => '0');
	channel_address_out <= wire_address_pres_reg_w_lg_w_q_range70w71w;
	channel_reconfig_done <= reconf_done_reg_out;
	clr_offset <= (is_offset_end AND en_mif_addr_cntr);
	default_max_limit_wire <= "1110";
	delay_mif_head_out <= delay_mif_head;
	delay_second_mif_head_out <= delay_second_mif_head;
	dprio_addr_index <= (wire_w_lg_w_lg_w_lg_w_lg_is_rx_pma515w516w518w519w OR wire_w_lg_w_lg_w_lg_is_rx_pma515w516w517w);
	dprio_addr_offset_cnt_out <= wire_dprio_addr_offset_cnt_q;
	dprio_addr_translated_offset <= (wire_add_sub6_w_lg_w_lg_result531w532w OR wire_w_lg_is_table_34529w);
	dprio_datain <= (wire_w_lg_w621w622w OR wire_w_lg_w_lg_is_tier_1613w614w);
	dprio_datain_64_67 <= (OTHERS => '0');
	dprio_datain_68_6B <= (OTHERS => '0');
	dprio_datain_preemp1t <= (OTHERS => '0');
	dprio_datain_vodctrl <= (OTHERS => '0');
	dprio_pulse <= ((dprio_pulse_reg XOR wire_dprio_busy) AND wire_dprio_w_lg_busy125w(0));
	dprio_wr_done <= wire_dprio_status_out(1);
	en_mif_addr_cntr <= ((read_state AND dprio_wr_done) OR wire_w_lg_w_lg_write_state384w385w(0));
	en_write_trigger <= '1';
	error <= error_reg;
	header_proc <= ((((delay_mif_head OR is_mif_header) OR delay_second_mif_head_out) OR is_second_mif_header) AND is_tier_1);
	idle_state <= (NOT state_mc_reg(0));
	invalid_eq_dcgain <= '0';
	is_ageb_table_7 <= ((wire_is_table_8_idx_ageb AND is_tier_1) AND is_rx_pcs);
	is_analog_control <= wire_reconf_mode_dec_eq(0);
	is_bonded_reconfig <= '0';
	is_central_pcs <= wire_reconf_mode_dec_eq(7);
	is_channel_reconfig <= wire_reconf_mode_dec_eq(1);
	is_end_mif <= end_mif_reg;
	is_illegal_reg_d <= (wire_w_lg_is_tier_218w(0) OR (wire_w_lg_w_lg_w25w26w27w(0) AND wire_w_lg_write_done19w(0)));
	is_illegal_reg_out <= is_illegal_reg;
	is_mif_header <= wire_is_special_address_aeb;
	is_mif_stage <= mif_stage;
	is_offset_end <= wire_dprio_addr_offset_cmpr_aeb;
	is_pma_mif_type <= (is_tx_pma OR is_rx_pma);
	is_protected_bit <= ((((((is_table_37 OR is_table_38) OR is_table_42) OR is_table_43) OR is_table_44) OR is_table_46) OR is_table_47);
	is_rcxpat_chnl_en_ch <= ((wire_is_rcxpat_chnl_en_ch_word_aeb AND is_tier_1) AND is_tx_pcs);
	is_rx_mif_type <= (is_rx_pcs OR is_rx_pma);
	is_rx_pcs <= (wire_mif_type_reg_w_lg_w_q_range495w496w(0) AND wire_w_lg_is_channel_reconfig491w(0));
	is_rx_pma <= (((wire_mif_type_reg_w_lg_w_q_range504w505w(0) AND wire_w_lg_is_rx_pcs498w(0)) AND wire_w_lg_is_tx_pma503w(0)) AND wire_w_lg_is_channel_reconfig491w(0));
	is_second_mif_header <= wire_is_second_mif_header_address_aeb;
	is_table_33 <= ((wire_is_table_33_idx_aeb AND is_tier_1) AND is_tx_pma);
	is_table_34 <= ((wire_is_table_34_idx_aeb AND is_tier_1) AND is_rx_pma);
	is_table_35 <= (wire_is_table_35_cmp_aeb AND is_tx_pma);
	is_table_37 <= ((wire_is_table_37_cmp_aeb AND is_tier_1) AND is_rx_pma);
	is_table_38 <= ((wire_is_table_38_cmp_aeb AND is_tier_1) AND is_rx_pma);
	is_table_42 <= ((wire_is_table_42_cmp_aeb AND is_tier_1) AND is_rx_pma);
	is_table_43 <= ((wire_is_table_43_cmp_aeb AND is_tier_1) AND is_rx_pma);
	is_table_44 <= ((wire_is_table_44_cmp_aeb AND is_tier_1) AND is_rx_pma);
	is_table_46 <= ((wire_is_table_46_cmp_aeb AND is_tier_1) AND is_rx_pma);
	is_table_47 <= ((wire_is_table_47_cmp_aeb AND is_tier_1) AND is_rx_pma);
	is_table_59 <= '0';
	is_table_61 <= '0';
	is_table_75 <= ((wire_is_table_75_idx_aeb AND is_tier_1) AND is_central_pcs);
	is_table_76 <= ((wire_is_table_76_idx_aeb AND is_tier_1) AND is_central_pcs);
	is_table_77 <= ((wire_is_table_77_idx_aeb AND is_tier_1) AND is_central_pcs);
	is_tier_1 <= (wire_reconf_mode_dec_eq(1) OR wire_reconf_mode_dec_eq(7));
	is_tier_2 <= wire_reconf_mode_dec_eq(2);
	is_tx_pcs <= wire_mif_type_reg_w_lg_w_q_range492w493w(0);
	is_tx_pma <= ((wire_mif_type_reg_w_lg_w_q_range499w500w(0) AND wire_w_lg_is_rx_pcs498w(0)) AND wire_w_lg_is_channel_reconfig491w(0));
	load_mif_header <= ((is_mif_header AND wire_w_lg_write_mif_word_done201w(0)) AND is_tier_1);
	merged_dprioin <= ( reconfig_data_reg(15 DOWNTO 12) & wire_w_lg_w_lg_w_lg_write_skip170w309w310w & wire_w319w & wire_w_lg_w_lg_w_lg_write_skip170w324w325w);
	mif_family_error <= ((NOT ((NOT reconfig_data_reg(7)) AND reconfig_data_reg(6))) AND is_second_mif_header);
	mif_reconfig_done <= ((wire_mif_type_reg_w_lg_w575w576w(0) AND wire_w_lg_is_central_pcs490w(0)) OR wire_w_lg_w_lg_is_central_pcs569w570w(0));
	mif_rx_only <= ((NOT mif_type_reg(1)) AND (NOT mif_type_reg(3)));
	mif_type_error <= ((((((NOT reconfig_data_reg(15)) AND (NOT reconfig_data_reg(14))) AND (NOT reconfig_data_reg(13))) AND (NOT reconfig_data_reg(12))) AND is_channel_reconfig) AND is_mif_header);
	offset_cancellation_reset <= '0';
	quad_address <= (OTHERS => '0');
	quad_address_out <= address_pres_reg(11 DOWNTO 3);
	rd_pulse <= ((((wire_w_lg_dprio_pulse146w(0) AND wire_w_lg_write_done19w(0)) AND wire_wr_rd_pulse_reg_w_lg_q128w(0)) AND wire_w_lg_is_illegal_reg_d163w(0)) AND wire_w_lg_write_state162w(0));
	read_address <= (OTHERS => '0');
	read_reconfig_addr <= (OTHERS => '0');
	read_state <= '0';
	reconf_done_reg_out <= reconfig_done_reg;
	reconfig_address_en <= (write_done OR idle_state);
	reconfig_address_out <= wire_mif_addr_cntr_w_lg_w_lg_q416w417w;
	reconfig_datain <= ((((((((((((wire_w_lg_is_table_33369w OR wire_w_lg_is_table_35368w) OR wire_w_lg_is_table_75367w) OR wire_w_lg_is_table_76366w) OR wire_w_lg_is_table_77365w) OR wire_w_lg_is_table_37364w) OR wire_w_lg_is_table_38363w) OR wire_w_lg_is_table_42362w) OR wire_w_lg_is_table_43361w) OR wire_w_lg_is_table_44360w) OR wire_w_lg_is_table_46359w) OR wire_w_lg_is_table_47358w) OR wire_w_lg_merged_dprioin357w);
	reconfig_reset_all <= reconfig_reset;
	reconfig_togxb <= ( wire_calibration_c3gxb_busy & wire_dprio_dprioload & wire_dprio_dpriodisable & wire_dprio_dprioin);
	reset_addr_done <= reconfig_reset_all;
	reset_reconf_addr <= '0';
	reset_system <= (wire_max_oper_limit_aeb AND wire_w_lg_idle_state31w(0));
	rx_pcs_max <= "10101";
	rx_pma_max <= "01100";
	rx_pma_minus_one <= "00001";
	rx_reconfig <= '1';
	s0_to_0 <= write_done;
	s0_to_1 <= (write_all_int AND idle_state);
	s0_to_2 <= '0';
	s2_to_0 <= '0';
	state_mc_reg_in(0) <= ((s0_to_2 OR s0_to_1) OR (((wire_w_lg_s2_to_010w(0) AND wire_w_lg_s0_to_19w(0)) AND wire_w_lg_s0_to_08w(0)) AND state_mc_reg(0)));
	table_33_data <= ( reconfig_data_reg(15 DOWNTO 0));
	table_34_addr <= "00110";
	table_35_data <= ( reconfig_data_reg(15 DOWNTO 0));
	table_37_data <= ( wire_w_lg_w_lg_w_lg_write_skip170w260w261w & dprio_dataout_reg(11 DOWNTO 3) & wire_w_lg_w_lg_w_lg_write_skip170w245w246w);
	table_38_data <= ( wire_w_lg_w_lg_w_lg_write_skip170w270w271w & dprio_dataout_reg(6 DOWNTO 5) & wire_w_lg_w_lg_w_lg_write_skip170w279w280w);
	table_42_data <= ( reconfig_data_reg(15 DOWNTO 0));
	table_43_data <= ( dprio_dataout_reg(15 DOWNTO 3) & wire_w_lg_w_lg_w_lg_write_skip170w245w246w);
	table_44_data <= ( wire_w_lg_w_lg_w_lg_write_skip170w290w291w);
	table_46_data <= ( dprio_dataout_reg(15 DOWNTO 10) & wire_w_lg_w_lg_w_lg_write_skip170w300w301w);
	table_47_data <= ( dprio_dataout_reg(15 DOWNTO 0));
	table_75_data <= ( wire_w_lg_w_lg_w_lg_write_skip170w212w213w & dprio_dataout_reg(14) & wire_w_lg_w_lg_w_lg_write_skip170w221w222w & dprio_dataout_reg(11) & wire_w_lg_w_lg_w_lg_write_skip170w229w230w);
	table_76_data <= ( dprio_dataout_reg(15) & wire_w_lg_w_lg_w_lg_write_skip170w237w238w & dprio_dataout_reg(5 DOWNTO 3) & wire_w_lg_w_lg_w_lg_write_skip170w245w246w);
	table_77_data <= ( dprio_dataout_reg(15 DOWNTO 14) & wire_w_lg_w_lg_w_lg_write_skip170w254w255w);
	tx_pcs_max <= "00011";
	tx_pma_max <= "00110";
	tx_reconfig <= '1';
	wr_pulse <= (((wire_w_lg_write_state181w(0) AND wire_w_lg_write_done19w(0)) AND (wire_wr_rd_pulse_reg_w_lg_q179w(0) OR (wire_w_lg_is_tier_1175w(0) AND ((wire_w_lg_w_lg_is_rcxpat_chnl_en_ch171w172w(0) AND wire_w_lg_bonded_skip169w(0)) AND wire_w_lg_is_protected_bit168w(0))))) AND wire_w_lg_is_illegal_reg_d163w(0));
	write_address <= ( "0" & address_pres_reg(2) & channel_address_out & "11" & "000000" & "0000");
	write_all_int <= (write_all AND en_write_trigger);
	write_done <= ((((wire_w_lg_w_lg_write_word_done633w634w(0) OR (wire_w_lg_w_lg_delay_mif_head_out630w631w(0) OR (reset_addr_done AND is_tier_1))) OR wire_w_lg_w_lg_dprio_pulse600w628w(0)) OR (is_illegal_reg_out AND write_state)) OR reset_system);
	write_happened <= wr_addr_inc_reg;
	write_mif_word_done <= (wire_w_lg_dprio_pulse600w(0) AND is_tier_1);
	write_reconfig_addr <= ( "0" & address_pres_reg(2) & wire_w_lg_w_channel_address_out_range669w670w & wire_w_lg_w_channel_address_out_range666w667w & wire_w_lg_is_pma_mif_type664w & wire_w_lg_w_lg_is_rx_mif_type661w662w & "00000" & dprio_addr_index(4 DOWNTO 1) & wire_w_lg_is_table_35648w);
	write_skip <= (((is_tx_pcs OR is_tx_pma) AND wire_w_lg_tx_reconfig21w(0)) OR ((is_rx_pcs OR is_rx_pma) AND wire_w_lg_rx_reconfig20w(0)));
	write_state <= state_mc_reg(0);
	write_word_64_67_data_valid <= '0';
	write_word_68_6B_data_valid <= '0';
	write_word_done <= '0';
	write_word_preemp1t_data_valid <= '0';
	write_word_vodctrl_data_valid <= '0';
	wire_w_cal_channel_address_range59w(0) <= cal_channel_address(0);
	wire_w_cal_channel_address_range53w(0) <= cal_channel_address(1);
	wire_w_cal_channel_address_range46w(0) <= cal_channel_address(2);
	wire_w_channel_address_range57w(0) <= channel_address(0);
	wire_w_channel_address_range50w(0) <= channel_address(1);
	wire_w_channel_address_out_range666w(0) <= channel_address_out(0);
	wire_w_channel_address_out_range669w(0) <= channel_address_out(1);
	wire_w_dprio_addr_index_range647w(0) <= dprio_addr_index(0);
	loop84 : FOR i IN 0 TO 15 GENERATE 
		wire_calibration_c3gxb_w_lg_w_lg_busy97w101w(i) <= wire_calibration_c3gxb_w_lg_busy97w(0) AND a2gr_dprio_addr(i);
	END GENERATE loop84;
	loop85 : FOR i IN 0 TO 15 GENERATE 
		wire_calibration_c3gxb_w_lg_w_lg_busy97w98w(i) <= wire_calibration_c3gxb_w_lg_busy97w(0) AND a2gr_dprio_data(i);
	END GENERATE loop85;
	wire_calibration_c3gxb_w_lg_w_lg_busy97w104w(0) <= wire_calibration_c3gxb_w_lg_busy97w(0) AND a2gr_dprio_rden;
	wire_calibration_c3gxb_w_lg_w_lg_busy97w107w(0) <= wire_calibration_c3gxb_w_lg_busy97w(0) AND a2gr_dprio_wren;
	wire_calibration_c3gxb_w_lg_w_lg_busy97w110w(0) <= wire_calibration_c3gxb_w_lg_busy97w(0) AND a2gr_dprio_wren_data;
	loop86 : FOR i IN 0 TO 15 GENERATE 
		wire_calibration_c3gxb_w_lg_busy102w(i) <= wire_calibration_c3gxb_busy AND cal_dprio_address(i);
	END GENERATE loop86;
	loop87 : FOR i IN 0 TO 15 GENERATE 
		wire_calibration_c3gxb_w_lg_busy99w(i) <= wire_calibration_c3gxb_busy AND wire_calibration_c3gxb_dprio_dataout(i);
	END GENERATE loop87;
	wire_calibration_c3gxb_w_lg_busy97w(0) <= NOT wire_calibration_c3gxb_busy;
	wire_calibration_c3gxb_reset <= wire_w_lg_offset_cancellation_reset82w(0);
	wire_w_lg_offset_cancellation_reset82w(0) <= offset_cancellation_reset OR reconfig_reset_all;
	calibration_c3gxb :  alt_cal_c3gxb
	  GENERIC MAP (
		CHANNEL_ADDRESS_WIDTH => 0,
		NUMBER_OF_CHANNELS => 1,
		SIM_MODEL_MODE => "FALSE"
	  )
	  PORT MAP ( 
		busy => wire_calibration_c3gxb_busy,
		clock => reconfig_clk,
		dprio_addr => wire_calibration_c3gxb_dprio_addr,
		dprio_busy => wire_dprio_busy,
		dprio_datain => wire_dprio_dataout,
		dprio_dataout => wire_calibration_c3gxb_dprio_dataout,
		dprio_rden => wire_calibration_c3gxb_dprio_rden,
		dprio_wren => wire_calibration_c3gxb_dprio_wren,
		quad_addr => wire_calibration_c3gxb_quad_addr,
		remap_addr => address_pres_reg,
		reset => wire_calibration_c3gxb_reset,
		retain_addr => wire_calibration_c3gxb_retain_addr,
		testbuses => cal_testbuses
	  );
	wire_dprio_w_lg_w_lg_w_status_out_range382w404w405w(0) <= wire_dprio_w_lg_w_status_out_range382w404w(0) AND reset_system;
	wire_dprio_w_lg_busy125w(0) <= NOT wire_dprio_busy;
	wire_dprio_w_lg_w_status_out_range382w404w(0) <= wire_dprio_w_status_out_range382w(0) OR wire_dprio_w_status_out_range403w(0);
	wire_dprio_address <= wire_calibration_c3gxb_w_lg_w_lg_busy102w103w;
	loop88 : FOR i IN 0 TO 15 GENERATE 
		wire_calibration_c3gxb_w_lg_w_lg_busy102w103w(i) <= wire_calibration_c3gxb_w_lg_busy102w(i) OR wire_calibration_c3gxb_w_lg_w_lg_busy97w101w(i);
	END GENERATE loop88;
	wire_dprio_datain <= wire_calibration_c3gxb_w_lg_w_lg_busy99w100w;
	loop89 : FOR i IN 0 TO 15 GENERATE 
		wire_calibration_c3gxb_w_lg_w_lg_busy99w100w(i) <= wire_calibration_c3gxb_w_lg_busy99w(i) OR wire_calibration_c3gxb_w_lg_w_lg_busy97w98w(i);
	END GENERATE loop89;
	wire_dprio_rden <= wire_calibration_c3gxb_w_lg_w_lg_busy105w106w(0);
	wire_calibration_c3gxb_w_lg_w_lg_busy105w106w(0) <= (wire_calibration_c3gxb_busy AND wire_calibration_c3gxb_dprio_rden) OR wire_calibration_c3gxb_w_lg_w_lg_busy97w104w(0);
	wire_dprio_wren <= wire_calibration_c3gxb_w_lg_w_lg_busy108w109w(0);
	wire_calibration_c3gxb_w_lg_w_lg_busy108w109w(0) <= (wire_calibration_c3gxb_busy AND wire_calibration_c3gxb_dprio_wren) OR wire_calibration_c3gxb_w_lg_w_lg_busy97w107w(0);
	wire_dprio_wren_data <= wire_calibration_c3gxb_w_lg_w_lg_busy111w112w(0);
	wire_calibration_c3gxb_w_lg_w_lg_busy111w112w(0) <= (wire_calibration_c3gxb_busy AND wire_calibration_c3gxb_retain_addr) OR wire_calibration_c3gxb_w_lg_w_lg_busy97w110w(0);
	wire_dprio_w_status_out_range382w(0) <= wire_dprio_status_out(1);
	wire_dprio_w_status_out_range403w(0) <= wire_dprio_status_out(3);
	dprio :  ALTGX_RECONFIG_CIV_alt_dprio_q9l
	  PORT MAP ( 
		address => wire_dprio_address,
		busy => wire_dprio_busy,
		datain => wire_dprio_datain,
		dataout => wire_dprio_dataout,
		dpclk => reconfig_clk,
		dpriodisable => wire_dprio_dpriodisable,
		dprioin => wire_dprio_dprioin,
		dprioload => wire_dprio_dprioload,
		dprioout => cal_dprioout_wire(0),
		quad_address => quad_address_out,
		rden => wire_dprio_rden,
		reset => reconfig_reset_all,
		status_out => wire_dprio_status_out,
		wren => wire_dprio_wren,
		wren_data => wire_dprio_wren_data
	  );
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN address_pres_reg <= (OTHERS => '0');
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN address_pres_reg <= ( wire_w_lg_w_lg_cal_busy41w42w & wire_w_lg_w_lg_cal_busy47w48w & wire_w_lg_w_lg_cal_busy54w55w & wire_w_lg_w_lg_cal_busy60w61w);
		END IF;
	END PROCESS;
	wire_address_pres_reg_w_lg_w_lg_w_q_range66w67w68w(0) <= wire_address_pres_reg_w_lg_w_q_range66w67w(0) AND wire_address_pres_reg_w_q_range64w(0);
	loop90 : FOR i IN 0 TO 1 GENERATE 
		wire_address_pres_reg_w_lg_w_q_range70w71w(i) <= wire_address_pres_reg_w_q_range70w(i) AND wire_address_pres_reg_w_lg_w_lg_w_lg_w_q_range66w67w68w69w(0);
	END GENERATE loop90;
	wire_address_pres_reg_w_lg_w_q_range66w67w(0) <= wire_address_pres_reg_w_q_range66w(0) AND wire_address_pres_reg_w_q_range65w(0);
	wire_address_pres_reg_w_lg_w_lg_w_lg_w_q_range66w67w68w69w(0) <= NOT wire_address_pres_reg_w_lg_w_lg_w_q_range66w67w68w(0);
	wire_address_pres_reg_w_q_range64w(0) <= address_pres_reg(0);
	wire_address_pres_reg_w_q_range70w <= address_pres_reg(1 DOWNTO 0);
	wire_address_pres_reg_w_q_range65w(0) <= address_pres_reg(1);
	wire_address_pres_reg_w_q_range66w(0) <= address_pres_reg(2);
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN delay_mif_head <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_delay_mif_head_ena = '1') THEN delay_mif_head <= (is_mif_header AND is_tier_1);
			END IF;
		END IF;
	END PROCESS;
	wire_delay_mif_head_ena <= (((wire_w_lg_write_state448w(0) AND wire_w_lg_write_mif_word_done201w(0)) AND wire_w_lg_reset_reconf_addr159w(0)) AND wire_w_lg_reset_system447w(0));
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN delay_second_mif_head <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_delay_second_mif_head_ena = '1') THEN delay_second_mif_head <= (is_second_mif_header AND wire_w_lg_write_done19w(0));
			END IF;
		END IF;
	END PROCESS;
	wire_delay_second_mif_head_ena <= (((wire_w_lg_write_state457w(0) AND wire_w_lg_reset_reconf_addr159w(0)) AND wire_w_lg_reset_system447w(0)) AND is_tier_1);
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN dprio_dataout_reg <= (OTHERS => '0');
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN dprio_dataout_reg <= wire_dprio_dataout;
		END IF;
	END PROCESS;
	wire_dprio_dataout_reg_w_q_range226w <= dprio_dataout_reg(10 DOWNTO 0);
	wire_dprio_dataout_reg_w_q_range264w <= dprio_dataout_reg(11 DOWNTO 3);
	wire_dprio_dataout_reg_w_q_range251w <= dprio_dataout_reg(13 DOWNTO 0);
	wire_dprio_dataout_reg_w_q_range218w <= dprio_dataout_reg(13 DOWNTO 12);
	wire_dprio_dataout_reg_w_q_range234w <= dprio_dataout_reg(14 DOWNTO 6);
	wire_dprio_dataout_reg_w_q_range288w <= dprio_dataout_reg(15 DOWNTO 0);
	wire_dprio_dataout_reg_w_q_range257w <= dprio_dataout_reg(15 DOWNTO 12);
	wire_dprio_dataout_reg_w_q_range209w(0) <= dprio_dataout_reg(15);
	wire_dprio_dataout_reg_w_q_range267w <= dprio_dataout_reg(15 DOWNTO 7);
	wire_dprio_dataout_reg_w_q_range242w <= dprio_dataout_reg(2 DOWNTO 0);
	wire_dprio_dataout_reg_w_q_range312w <= dprio_dataout_reg(2 DOWNTO 1);
	wire_dprio_dataout_reg_w_q_range276w <= dprio_dataout_reg(4 DOWNTO 0);
	wire_dprio_dataout_reg_w_q_range297w <= dprio_dataout_reg(9 DOWNTO 0);
	wire_dprio_dataout_reg_w_q_range321w(0) <= dprio_dataout_reg(0);
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN dprio_pulse_reg <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_dprio_pulse_reg_ena = '1') THEN dprio_pulse_reg <= wire_dprio_busy;
			END IF;
		END IF;
	END PROCESS;
	wire_dprio_pulse_reg_ena <= (read_state OR write_state);
	PROCESS (reconfig_clk)
	BEGIN
		IF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (is_tier_1 = '1') THEN end_mif_reg <= mif_reconfig_done;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN error_reg <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN error_reg <= (is_illegal_reg OR reset_system);
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN is_illegal_reg <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN is_illegal_reg <= (((wire_w_lg_is_illegal_reg_d35w(0) AND wire_w_lg_is_illegal_reg_out34w(0)) OR (is_illegal_reg_out AND write_done)) OR reset_system);
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, wire_mif_central_pcs_error_reg_clrn)
	BEGIN
		IF (wire_mif_central_pcs_error_reg_clrn = '0') THEN mif_central_pcs_error_reg <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (delay_second_mif_head_out = '1') THEN mif_central_pcs_error_reg <= ((NOT reconfig_data_reg(15)) AND is_central_pcs);
			END IF;
		END IF;
	END PROCESS;
	wire_mif_central_pcs_error_reg_clrn <= (NOT (reset_addr_done OR is_illegal_reg_out));
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN mif_stage <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (is_tier_1 = '1') THEN 
				IF (wire_mif_stage_sclr = '1') THEN mif_stage <= '0';
				ELSE mif_stage <= ((wire_mif_stage_w_lg_q194w(0) AND wire_w_lg_is_mif_header190w(0)) OR wire_w_lg_w_lg_w_lg_w_lg_is_mif_header190w191w192w193w(0));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	wire_mif_stage_sclr <= ((reset_system OR is_illegal_reg_out) OR mif_reconfig_done);
	wire_mif_stage_w_lg_q194w(0) <= NOT mif_stage;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN mif_type_reg(0) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_mif_type_reg_ena(0) = '1') THEN 
				IF (wire_mif_type_reg_sclr(0) = '1') THEN mif_type_reg(0) <= '0';
				ELSE mif_type_reg(0) <= wire_mif_type_reg_d(0);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN mif_type_reg(1) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_mif_type_reg_ena(1) = '1') THEN 
				IF (wire_mif_type_reg_sclr(1) = '1') THEN mif_type_reg(1) <= '0';
				ELSE mif_type_reg(1) <= wire_mif_type_reg_d(1);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN mif_type_reg(2) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_mif_type_reg_ena(2) = '1') THEN 
				IF (wire_mif_type_reg_sclr(2) = '1') THEN mif_type_reg(2) <= '0';
				ELSE mif_type_reg(2) <= wire_mif_type_reg_d(2);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN mif_type_reg(3) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_mif_type_reg_ena(3) = '1') THEN 
				IF (wire_mif_type_reg_sclr(3) = '1') THEN mif_type_reg(3) <= '0';
				ELSE mif_type_reg(3) <= wire_mif_type_reg_d(3);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	wire_mif_type_reg_d <= wire_reconfig_data_reg_w_lg_w_lg_w_lg_w_q_range259w476w477w478w;
	loop91 : FOR i IN 0 TO 3 GENERATE
		wire_mif_type_reg_ena(i) <= wire_w_lg_load_mif_header473w(0);
	END GENERATE loop91;
	wire_mif_type_reg_sclr <= ( wire_w_lg_w_lg_w_lg_load_mif_header479w480w481w & wire_w_lg_w_lg_w_lg_load_mif_header479w480w484w & wire_w_lg_w_lg_w_lg_load_mif_header479w480w486w & wire_w_lg_w_lg_w_lg_load_mif_header479w480w488w);
	wire_mif_type_reg_w_lg_w575w576w(0) <= wire_mif_type_reg_w575w(0) AND write_done;
	wire_mif_type_reg_w_lg_w_lg_w_lg_w_lg_w_q_range492w571w572w573w574w(0) <= wire_mif_type_reg_w_lg_w_lg_w_lg_w_q_range492w571w572w573w(0) AND is_channel_reconfig;
	wire_mif_type_reg_w_lg_w_q_range504w505w(0) <= wire_mif_type_reg_w_q_range504w(0) AND wire_w_lg_is_tx_pcs494w(0);
	wire_mif_type_reg_w_lg_w_q_range499w500w(0) <= wire_mif_type_reg_w_q_range499w(0) AND wire_w_lg_is_tx_pcs494w(0);
	wire_mif_type_reg_w_lg_w_q_range495w496w(0) <= wire_mif_type_reg_w_q_range495w(0) AND wire_w_lg_is_tx_pcs494w(0);
	wire_mif_type_reg_w_lg_w_q_range492w493w(0) <= wire_mif_type_reg_w_q_range492w(0) AND wire_w_lg_is_channel_reconfig491w(0);
	wire_mif_type_reg_w575w(0) <= NOT wire_mif_type_reg_w_lg_w_lg_w_lg_w_lg_w_q_range492w571w572w573w574w(0);
	wire_mif_type_reg_w_lg_w_lg_w_lg_w_q_range492w571w572w573w(0) <= wire_mif_type_reg_w_lg_w_lg_w_q_range492w571w572w(0) OR wire_mif_type_reg_w_q_range504w(0);
	wire_mif_type_reg_w_lg_w_lg_w_q_range492w571w572w(0) <= wire_mif_type_reg_w_lg_w_q_range492w571w(0) OR wire_mif_type_reg_w_q_range499w(0);
	wire_mif_type_reg_w_lg_w_q_range492w571w(0) <= wire_mif_type_reg_w_q_range492w(0) OR wire_mif_type_reg_w_q_range495w(0);
	wire_mif_type_reg_w_q_range504w(0) <= mif_type_reg(0);
	wire_mif_type_reg_w_q_range499w(0) <= mif_type_reg(1);
	wire_mif_type_reg_w_q_range495w(0) <= mif_type_reg(2);
	wire_mif_type_reg_w_q_range492w(0) <= mif_type_reg(3);
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN reconf_mode_sel_reg(0) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_reconf_mode_sel_reg_ena(0) = '1') THEN reconf_mode_sel_reg(0) <= reconfig_mode_sel(0);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN reconf_mode_sel_reg(1) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_reconf_mode_sel_reg_ena(1) = '1') THEN reconf_mode_sel_reg(1) <= reconfig_mode_sel(1);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN reconf_mode_sel_reg(2) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_reconf_mode_sel_reg_ena(2) = '1') THEN reconf_mode_sel_reg(2) <= reconfig_mode_sel(2);
			END IF;
		END IF;
	END PROCESS;
	loop92 : FOR i IN 0 TO 2 GENERATE
		wire_reconf_mode_sel_reg_ena(i) <= wire_w_lg_idle_state200w(0);
	END GENERATE loop92;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN reconfig_data_reg(0) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_reconfig_data_reg_ena(0) = '1') THEN reconfig_data_reg(0) <= reconfig_data(0);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN reconfig_data_reg(1) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_reconfig_data_reg_ena(1) = '1') THEN reconfig_data_reg(1) <= reconfig_data(1);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN reconfig_data_reg(2) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_reconfig_data_reg_ena(2) = '1') THEN reconfig_data_reg(2) <= reconfig_data(2);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN reconfig_data_reg(3) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_reconfig_data_reg_ena(3) = '1') THEN reconfig_data_reg(3) <= reconfig_data(3);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN reconfig_data_reg(4) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_reconfig_data_reg_ena(4) = '1') THEN reconfig_data_reg(4) <= reconfig_data(4);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN reconfig_data_reg(5) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_reconfig_data_reg_ena(5) = '1') THEN reconfig_data_reg(5) <= reconfig_data(5);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN reconfig_data_reg(6) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_reconfig_data_reg_ena(6) = '1') THEN reconfig_data_reg(6) <= reconfig_data(6);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN reconfig_data_reg(7) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_reconfig_data_reg_ena(7) = '1') THEN reconfig_data_reg(7) <= reconfig_data(7);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN reconfig_data_reg(8) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_reconfig_data_reg_ena(8) = '1') THEN reconfig_data_reg(8) <= reconfig_data(8);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN reconfig_data_reg(9) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_reconfig_data_reg_ena(9) = '1') THEN reconfig_data_reg(9) <= reconfig_data(9);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN reconfig_data_reg(10) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_reconfig_data_reg_ena(10) = '1') THEN reconfig_data_reg(10) <= reconfig_data(10);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN reconfig_data_reg(11) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_reconfig_data_reg_ena(11) = '1') THEN reconfig_data_reg(11) <= reconfig_data(11);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN reconfig_data_reg(12) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_reconfig_data_reg_ena(12) = '1') THEN reconfig_data_reg(12) <= reconfig_data(12);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN reconfig_data_reg(13) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_reconfig_data_reg_ena(13) = '1') THEN reconfig_data_reg(13) <= reconfig_data(13);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN reconfig_data_reg(14) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_reconfig_data_reg_ena(14) = '1') THEN reconfig_data_reg(14) <= reconfig_data(14);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN reconfig_data_reg(15) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_reconfig_data_reg_ena(15) = '1') THEN reconfig_data_reg(15) <= reconfig_data(15);
			END IF;
		END IF;
	END PROCESS;
	loop93 : FOR i IN 0 TO 15 GENERATE
		wire_reconfig_data_reg_ena(i) <= wire_w_lg_idle_state327w(0);
	END GENERATE loop93;
	loop94 : FOR i IN 0 TO 3 GENERATE 
		wire_reconfig_data_reg_w_lg_w_lg_w_q_range259w476w477w(i) <= wire_reconfig_data_reg_w_lg_w_q_range259w476w(i) AND wire_w_lg_clr_offset475w(0);
	END GENERATE loop94;
	loop95 : FOR i IN 0 TO 3 GENERATE 
		wire_reconfig_data_reg_w_lg_w_q_range259w476w(i) <= wire_reconfig_data_reg_w_q_range259w(i) AND load_mif_header;
	END GENERATE loop95;
	loop96 : FOR i IN 0 TO 3 GENERATE 
		wire_reconfig_data_reg_w_lg_w_lg_w_lg_w_q_range259w476w477w478w(i) <= wire_reconfig_data_reg_w_lg_w_lg_w_q_range259w476w477w(i) OR wire_w_lg_clr_offset474w(i);
	END GENERATE loop96;
	wire_reconfig_data_reg_w_q_range323w(0) <= reconfig_data_reg(0);
	wire_reconfig_data_reg_w_q_range228w <= reconfig_data_reg(10 DOWNTO 0);
	wire_reconfig_data_reg_w_q_range308w <= reconfig_data_reg(11 DOWNTO 3);
	wire_reconfig_data_reg_w_q_range253w <= reconfig_data_reg(13 DOWNTO 0);
	wire_reconfig_data_reg_w_q_range220w <= reconfig_data_reg(13 DOWNTO 12);
	wire_reconfig_data_reg_w_q_range236w <= reconfig_data_reg(14 DOWNTO 6);
	wire_reconfig_data_reg_w_q_range204w <= reconfig_data_reg(15 DOWNTO 0);
	wire_reconfig_data_reg_w_q_range259w <= reconfig_data_reg(15 DOWNTO 12);
	wire_reconfig_data_reg_w_q_range211w(0) <= reconfig_data_reg(15);
	wire_reconfig_data_reg_w_q_range269w <= reconfig_data_reg(15 DOWNTO 7);
	wire_reconfig_data_reg_w_q_range244w <= reconfig_data_reg(2 DOWNTO 0);
	wire_reconfig_data_reg_w_q_range314w <= reconfig_data_reg(2 DOWNTO 1);
	wire_reconfig_data_reg_w_q_range278w <= reconfig_data_reg(4 DOWNTO 0);
	wire_reconfig_data_reg_w_q_range299w <= reconfig_data_reg(9 DOWNTO 0);
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN reconfig_done_reg <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_reconfig_done_reg_ena = '1') THEN 
				IF (reset_system = '1') THEN reconfig_done_reg <= '0';
				ELSE reconfig_done_reg <= (((mif_reconfig_done AND is_tier_1) AND wire_reconfig_done_reg_w_lg_q469w(0)) OR wire_reconfig_done_reg_w_lg_q468w(0));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	wire_reconfig_done_reg_ena <= (is_mif_stage OR (idle_state AND wire_w_lg_is_mif_stage461w(0)));
	wire_reconfig_done_reg_w_lg_q468w(0) <= reconfig_done_reg AND wire_w_lg_w_lg_w_lg_is_mif_header465w466w467w(0);
	wire_reconfig_done_reg_w_lg_q469w(0) <= NOT reconfig_done_reg;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN state_mc_reg <= (OTHERS => '0');
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN state_mc_reg <= state_mc_reg_in;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN wr_addr_inc_reg <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN wr_addr_inc_reg <= (wr_pulse OR ((wire_w_lg_wr_pulse74w(0) AND wire_w_lg_rd_pulse73w(0)) AND wr_addr_inc_reg));
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN wr_rd_pulse_reg <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_wr_rd_pulse_reg_ena = '1') THEN 
				IF (wire_wr_rd_pulse_reg_sclr = '1') THEN wr_rd_pulse_reg <= '0';
				ELSE wr_rd_pulse_reg <= wire_wr_rd_pulse_reg_w_lg_q128w(0);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	wire_wr_rd_pulse_reg_ena <= (((((wire_w_lg_dprio_pulse146w(0) AND wire_w_lg_delay_mif_head_out145w(0)) OR (wire_w_lg_dprio_pulse139w(0) AND wire_w_lg_read_state130w(0))) OR (is_tier_1 AND mif_reconfig_done)) OR reset_addr_done) OR is_illegal_reg_out);
	wire_wr_rd_pulse_reg_sclr <= (((reset_system OR (is_tier_1 AND mif_reconfig_done)) OR reset_addr_done) OR is_illegal_reg_out);
	wire_wr_rd_pulse_reg_w_lg_q179w(0) <= wr_rd_pulse_reg AND wire_w_lg_w_lg_is_tier_1137w178w(0);
	wire_wr_rd_pulse_reg_w_lg_q128w(0) <= NOT wr_rd_pulse_reg;
	PROCESS (reconfig_clk, wire_wren_data_reg_clrn)
	BEGIN
		IF (wire_wren_data_reg_clrn = '0') THEN wren_data_reg <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_wren_data_reg_ena = '1') THEN wren_data_reg <= rd_pulse;
			END IF;
		END IF;
	END PROCESS;
	wire_wren_data_reg_clrn <= (NOT (write_done OR reconfig_reset_all));
	wire_wren_data_reg_ena <= (rd_pulse AND is_tier_1);
	wire_wren_data_reg_w_lg_q608w(0) <= NOT wren_data_reg;
	loop97 : FOR i IN 0 TO 4 GENERATE 
		wire_add_sub6_w_lg_w_lg_result531w532w(i) <= wire_add_sub6_w_lg_result531w(i) AND wire_w_lg_is_table_34530w(0);
	END GENERATE loop97;
	loop98 : FOR i IN 0 TO 4 GENERATE 
		wire_add_sub6_w_lg_result531w(i) <= wire_add_sub6_result(i) AND wire_w_lg_w_lg_is_rx_pma515w516w(0);
	END GENERATE loop98;
	add_sub6 :  lpm_add_sub
	  GENERIC MAP (
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 5
	  )
	  PORT MAP ( 
		add_sub => add_sub_sel,
		dataa => wire_dprio_addr_offset_cnt_q,
		datab => add_sub_datab,
		result => wire_add_sub6_result
	  );
	wire_dprio_addr_offset_cmpr_datab <= wire_w_lg_w_lg_w_lg_is_central_pcs490w543w544w;
	loop99 : FOR i IN 0 TO 4 GENERATE 
		wire_w_lg_w_lg_w_lg_is_central_pcs490w543w544w(i) <= wire_w_lg_w_lg_is_central_pcs490w543w(i) OR wire_w_lg_is_central_pcs542w(i);
	END GENERATE loop99;
	dprio_addr_offset_cmpr :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 5
	  )
	  PORT MAP ( 
		aeb => wire_dprio_addr_offset_cmpr_aeb,
		dataa => wire_dprio_addr_offset_cnt_q,
		datab => wire_dprio_addr_offset_cmpr_datab
	  );
	wire_is_rcxpat_chnl_en_ch_word_datab <= "00001";
	is_rcxpat_chnl_en_ch_word :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 5
	  )
	  PORT MAP ( 
		aeb => wire_is_rcxpat_chnl_en_ch_word_aeb,
		dataa => dprio_addr_offset_cnt_out,
		datab => wire_is_rcxpat_chnl_en_ch_word_datab
	  );
	wire_is_second_mif_header_address_datab <= "000001";
	is_second_mif_header_address :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 6
	  )
	  PORT MAP ( 
		aeb => wire_is_second_mif_header_address_aeb,
		dataa => wire_mif_addr_cntr_q,
		datab => wire_is_second_mif_header_address_datab
	  );
	wire_is_special_address_datab <= (OTHERS => '0');
	is_special_address :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 6
	  )
	  PORT MAP ( 
		aeb => wire_is_special_address_aeb,
		dataa => wire_mif_addr_cntr_q,
		datab => wire_is_special_address_datab
	  );
	wire_is_table_33_idx_datab <= "00101";
	is_table_33_idx :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 5
	  )
	  PORT MAP ( 
		aeb => wire_is_table_33_idx_aeb,
		dataa => dprio_addr_offset_cnt_out,
		datab => wire_is_table_33_idx_datab
	  );
	wire_is_table_34_idx_datab <= (OTHERS => '0');
	is_table_34_idx :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 5
	  )
	  PORT MAP ( 
		aeb => wire_is_table_34_idx_aeb,
		dataa => dprio_addr_offset_cnt_out,
		datab => wire_is_table_34_idx_datab
	  );
	wire_is_table_35_cmp_datab <= "00110";
	is_table_35_cmp :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 5
	  )
	  PORT MAP ( 
		aeb => wire_is_table_35_cmp_aeb,
		dataa => dprio_addr_offset_cnt_out,
		datab => wire_is_table_35_cmp_datab
	  );
	wire_is_table_37_cmp_datab <= "00010";
	is_table_37_cmp :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 5
	  )
	  PORT MAP ( 
		aeb => wire_is_table_37_cmp_aeb,
		dataa => dprio_addr_offset_cnt_out,
		datab => wire_is_table_37_cmp_datab
	  );
	wire_is_table_38_cmp_datab <= "00011";
	is_table_38_cmp :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 5
	  )
	  PORT MAP ( 
		aeb => wire_is_table_38_cmp_aeb,
		dataa => dprio_addr_offset_cnt_out,
		datab => wire_is_table_38_cmp_datab
	  );
	wire_is_table_42_cmp_datab <= "00111";
	is_table_42_cmp :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 5
	  )
	  PORT MAP ( 
		aeb => wire_is_table_42_cmp_aeb,
		dataa => dprio_addr_offset_cnt_out,
		datab => wire_is_table_42_cmp_datab
	  );
	wire_is_table_43_cmp_datab <= "01000";
	is_table_43_cmp :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 5
	  )
	  PORT MAP ( 
		aeb => wire_is_table_43_cmp_aeb,
		dataa => dprio_addr_offset_cnt_out,
		datab => wire_is_table_43_cmp_datab
	  );
	wire_is_table_44_cmp_datab <= "01001";
	is_table_44_cmp :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 5
	  )
	  PORT MAP ( 
		aeb => wire_is_table_44_cmp_aeb,
		dataa => dprio_addr_offset_cnt_out,
		datab => wire_is_table_44_cmp_datab
	  );
	wire_is_table_46_cmp_datab <= "01011";
	is_table_46_cmp :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 5
	  )
	  PORT MAP ( 
		aeb => wire_is_table_46_cmp_aeb,
		dataa => dprio_addr_offset_cnt_out,
		datab => wire_is_table_46_cmp_datab
	  );
	wire_is_table_47_cmp_datab <= "01100";
	is_table_47_cmp :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 5
	  )
	  PORT MAP ( 
		aeb => wire_is_table_47_cmp_aeb,
		dataa => dprio_addr_offset_cnt_out,
		datab => wire_is_table_47_cmp_datab
	  );
	wire_is_table_75_idx_datab <= "00001";
	is_table_75_idx :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 5
	  )
	  PORT MAP ( 
		aeb => wire_is_table_75_idx_aeb,
		dataa => dprio_addr_offset_cnt_out,
		datab => wire_is_table_75_idx_datab
	  );
	wire_is_table_76_idx_datab <= "00010";
	is_table_76_idx :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 5
	  )
	  PORT MAP ( 
		aeb => wire_is_table_76_idx_aeb,
		dataa => dprio_addr_offset_cnt_out,
		datab => wire_is_table_76_idx_datab
	  );
	wire_is_table_77_idx_datab <= "00011";
	is_table_77_idx :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 5
	  )
	  PORT MAP ( 
		aeb => wire_is_table_77_idx_aeb,
		dataa => dprio_addr_offset_cnt_out,
		datab => wire_is_table_77_idx_datab
	  );
	wire_is_table_8_idx_datab <= "00010";
	is_table_8_idx :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 5
	  )
	  PORT MAP ( 
		ageb => wire_is_table_8_idx_ageb,
		dataa => dprio_addr_offset_cnt_out,
		datab => wire_is_table_8_idx_datab
	  );
	max_oper_limit :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 4
	  )
	  PORT MAP ( 
		aeb => wire_max_oper_limit_aeb,
		dataa => wire_oper_count_q,
		datab => default_max_limit_wire
	  );
	wire_dprio_addr_offset_cnt_data <= (OTHERS => '0');
	wire_dprio_addr_offset_cnt_sclr <= wire_w_lg_w_lg_w_lg_w_lg_clr_offset511w512w513w514w(0);
	wire_w_lg_w_lg_w_lg_w_lg_clr_offset511w512w513w514w(0) <= (((clr_offset OR is_mif_header) OR reset_addr_done) OR is_illegal_reg_out) OR mif_reconfig_done;
	dprio_addr_offset_cnt :  lpm_counter
	  GENERIC MAP (
		lpm_port_updown => "PORT_UNUSED",
		lpm_width => 5
	  )
	  PORT MAP ( 
		clock => reconfig_clk,
		cnt_en => en_mif_addr_cntr,
		data => wire_dprio_addr_offset_cnt_data,
		q => wire_dprio_addr_offset_cnt_q,
		sclr => wire_dprio_addr_offset_cnt_sclr
	  );
	loop100 : FOR i IN 0 TO 5 GENERATE 
		wire_mif_addr_cntr_w_lg_w_lg_q416w417w(i) <= wire_mif_addr_cntr_w_lg_q416w(i) AND is_tier_1;
	END GENERATE loop100;
	loop101 : FOR i IN 0 TO 5 GENERATE 
		wire_mif_addr_cntr_w_lg_q416w(i) <= wire_mif_addr_cntr_q(i) AND wire_w_lg_w_lg_mif_reconfig_done389w415w(0);
	END GENERATE loop101;
	wire_mif_addr_cntr_cnt_en <= wire_w_lg_w_lg_en_mif_addr_cntr397w398w(0);
	wire_w_lg_w_lg_en_mif_addr_cntr397w398w(0) <= (en_mif_addr_cntr OR ((((((is_mif_header AND write_state) OR (is_second_mif_header AND write_state)) AND wire_w_lg_write_done19w(0)) AND wire_w_lg_mif_reconfig_done389w(0)) AND wire_w_lg_reconf_done_reg_out388w(0)) AND wire_w_lg_dprio_pulse146w(0))) AND is_tier_1;
	wire_mif_addr_cntr_data <= wire_w_lg_is_central_pcs402w;
	wire_mif_addr_cntr_sclr <= wire_w_lg_w412w413w(0);
	wire_w_lg_w412w413w(0) <= ((((reset_reconf_addr OR is_end_mif) AND (NOT ((is_mif_header OR is_second_mif_header) AND write_state))) OR wire_dprio_w_lg_w_lg_w_status_out_range382w404w405w(0)) OR is_illegal_reg_out) OR reconfig_reset_all;
	wire_mif_addr_cntr_sload <= wire_w_lg_w_lg_w_lg_is_second_mif_header399w400w401w(0);
	wire_w_lg_w_lg_w_lg_is_second_mif_header399w400w401w(0) <= ((is_second_mif_header AND wire_w_lg_write_done19w(0)) AND write_state) AND is_central_pcs;
	mif_addr_cntr :  lpm_counter
	  GENERIC MAP (
		lpm_modulus => 50,
		lpm_port_updown => "PORT_UNUSED",
		lpm_width => 6
	  )
	  PORT MAP ( 
		clock => reconfig_clk,
		cnt_en => wire_mif_addr_cntr_cnt_en,
		data => wire_mif_addr_cntr_data,
		q => wire_mif_addr_cntr_q,
		sclr => wire_mif_addr_cntr_sclr,
		sload => wire_mif_addr_cntr_sload
	  );
	wire_oper_count_sclr <= wire_w_lg_idle_state30w(0);
	wire_w_lg_idle_state30w(0) <= idle_state OR reconfig_reset_all;
	oper_count :  lpm_counter
	  GENERIC MAP (
		lpm_port_updown => "PORT_UNUSED",
		lpm_width => 4
	  )
	  PORT MAP ( 
		clock => reconfig_clk,
		cnt_en => dprio_pulse,
		q => wire_oper_count_q,
		sclr => wire_oper_count_sclr
	  );
	wire_reconf_mode_dec_enable <= wire_w_lg_w_lg_idle_state31w199w(0);
	wire_w_lg_w_lg_idle_state31w199w(0) <= wire_w_lg_idle_state31w(0) OR mif_stage;
	reconf_mode_dec :  lpm_decode
	  GENERIC MAP (
		LPM_DECODES => 8,
		LPM_WIDTH => 3
	  )
	  PORT MAP ( 
		data => reconf_mode_sel_reg,
		enable => wire_reconf_mode_dec_enable,
		eq => wire_reconf_mode_dec_eq
	  );
	wire_central_pcs_first_word_mux_data <= ( "100101" & "001111" & "110000" & "001101" & "010110" & "001001");
	wire_central_pcs_first_word_mux_sel <= ( mif_rx_only & mif_type_reg(3) & wire_w_lg_w_lg_w_lg_mif_rx_only562w563w564w);
	central_pcs_first_word_mux :  ALTGX_RECONFIG_CIV_mux_cda
	  PORT MAP ( 
		data => wire_central_pcs_first_word_mux_data,
		result => wire_central_pcs_first_word_mux_result,
		sel => wire_central_pcs_first_word_mux_sel
	  );
	wire_max_word_per_mif_type_data <= ( rx_pma_max & tx_pma_max & rx_pcs_max & tx_pcs_max);
	wire_max_word_per_mif_type_sel <= ( is_pma_mif_type & is_rx_mif_type);
	max_word_per_mif_type :  ALTGX_RECONFIG_CIV_mux_8da
	  PORT MAP ( 
		data => wire_max_word_per_mif_type_data,
		result => wire_max_word_per_mif_type_result,
		sel => wire_max_word_per_mif_type_sel
	  );

 END RTL; --ALTGX_RECONFIG_CIV_alt_c3gxb_reconfig_osa1
--VALID FILE


LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY ALTGX_RECONFIG_CIV IS
	PORT
	(
		reconfig_clk		: IN STD_LOGIC ;
		reconfig_data		: IN STD_LOGIC_VECTOR (15 DOWNTO 0);
		reconfig_fromgxb		: IN STD_LOGIC_VECTOR (4 DOWNTO 0);
		reconfig_reset		: IN STD_LOGIC ;
		write_all		: IN STD_LOGIC ;
		busy		: OUT STD_LOGIC ;
		channel_reconfig_done		: OUT STD_LOGIC ;
		error		: OUT STD_LOGIC ;
		reconfig_address_en		: OUT STD_LOGIC ;
		reconfig_address_out		: OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
		reconfig_togxb		: OUT STD_LOGIC_VECTOR (3 DOWNTO 0)
	);
END ALTGX_RECONFIG_CIV;


ARCHITECTURE RTL OF altgx_reconfig_civ IS

	ATTRIBUTE synthesis_clearbox: natural;
	ATTRIBUTE synthesis_clearbox OF RTL: ARCHITECTURE IS 2;
	ATTRIBUTE clearbox_macroname: string;
	ATTRIBUTE clearbox_macroname OF RTL: ARCHITECTURE IS "alt_c3gxb_reconfig";
	ATTRIBUTE clearbox_defparam: string;
	ATTRIBUTE clearbox_defparam OF RTL: ARCHITECTURE IS "cbx_blackbox_list=-lpm_mux;enable_illegal_mode_check=TRUE;enable_self_recovery=TRUE;intended_device_family=Cyclone IV GX;mif_address_width=6;number_of_channels=1;number_of_reconfig_ports=1;enable_buf_cal=true;reconfig_fromgxb_width=5;reconfig_togxb_width=4;";
	SIGNAL sub_wire0	: STD_LOGIC ;
	SIGNAL sub_wire1	: STD_LOGIC ;
	SIGNAL sub_wire2	: STD_LOGIC ;
	SIGNAL sub_wire3	: STD_LOGIC ;
	SIGNAL sub_wire4	: STD_LOGIC_VECTOR (5 DOWNTO 0);
	SIGNAL sub_wire5	: STD_LOGIC_VECTOR (3 DOWNTO 0);
	SIGNAL sub_wire6_bv	: BIT_VECTOR (0 DOWNTO 0);
	SIGNAL sub_wire6	: STD_LOGIC_VECTOR (0 DOWNTO 0);
	SIGNAL sub_wire7	: STD_LOGIC_VECTOR (2 DOWNTO 0);
	SIGNAL sub_wire8_bv	: BIT_VECTOR (0 DOWNTO 0);
	SIGNAL sub_wire8	: STD_LOGIC_VECTOR (0 DOWNTO 0);



	COMPONENT ALTGX_RECONFIG_CIV_alt_c3gxb_reconfig_osa1
	PORT (
			reconfig_clk	: IN STD_LOGIC ;
			reconfig_data	: IN STD_LOGIC_VECTOR (15 DOWNTO 0);
			reconfig_fromgxb	: IN STD_LOGIC_VECTOR (4 DOWNTO 0);
			reconfig_mode_sel	: IN STD_LOGIC_VECTOR (2 DOWNTO 0);
			reconfig_reset	: IN STD_LOGIC ;
			write_all	: IN STD_LOGIC ;
			busy	: OUT STD_LOGIC ;
			channel_reconfig_done	: OUT STD_LOGIC ;
			error	: OUT STD_LOGIC ;
			reconfig_address_en	: OUT STD_LOGIC ;
			reconfig_address_out	: OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
			reconfig_togxb	: OUT STD_LOGIC_VECTOR (3 DOWNTO 0)
	);
	END COMPONENT;

BEGIN
	sub_wire6_bv(0 DOWNTO 0) <= "0";
	sub_wire6    <= NOT(To_stdlogicvector(sub_wire6_bv));
	sub_wire8_bv(0 DOWNTO 0) <= "0";
	sub_wire8    <= To_stdlogicvector(sub_wire8_bv);
	busy    <= sub_wire0;
	channel_reconfig_done    <= sub_wire1;
	error    <= sub_wire2;
	reconfig_address_en    <= sub_wire3;
	reconfig_address_out    <= sub_wire4(5 DOWNTO 0);
	reconfig_togxb    <= sub_wire5(3 DOWNTO 0);
	sub_wire7    <= sub_wire8(0 DOWNTO 0) & sub_wire8(0 DOWNTO 0) & sub_wire6(0 DOWNTO 0);

	ALTGX_RECONFIG_CIV_alt_c3gxb_reconfig_osa1_component : ALTGX_RECONFIG_CIV_alt_c3gxb_reconfig_osa1
	PORT MAP (
		reconfig_clk => reconfig_clk,
		reconfig_data => reconfig_data,
		reconfig_fromgxb => reconfig_fromgxb,
		reconfig_mode_sel => sub_wire7,
		reconfig_reset => reconfig_reset,
		write_all => write_all,
		busy => sub_wire0,
		channel_reconfig_done => sub_wire1,
		error => sub_wire2,
		reconfig_address_en => sub_wire3,
		reconfig_address_out => sub_wire4,
		reconfig_togxb => sub_wire5
	);



END RTL;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: ADCE NUMERIC "0"
-- Retrieval info: PRIVATE: CMU_PLL NUMERIC "0"
-- Retrieval info: PRIVATE: DATA_RATE NUMERIC "0"
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone IV GX"
-- Retrieval info: PRIVATE: PMA NUMERIC "0"
-- Retrieval info: PRIVATE: PROTO_SWITCH NUMERIC "1"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: CONSTANT: CBX_BLACKBOX_LIST STRING "-lpm_mux"
-- Retrieval info: CONSTANT: ENABLE_ILLEGAL_MODE_CHECK STRING "TRUE"
-- Retrieval info: CONSTANT: ENABLE_SELF_RECOVERY STRING "TRUE"
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone IV GX"
-- Retrieval info: CONSTANT: MIF_ADDRESS_WIDTH NUMERIC "6"
-- Retrieval info: CONSTANT: NUMBER_OF_CHANNELS NUMERIC "1"
-- Retrieval info: CONSTANT: NUMBER_OF_RECONFIG_PORTS NUMERIC "1"
-- Retrieval info: CONSTANT: enable_buf_cal STRING "true"
-- Retrieval info: CONSTANT: reconfig_fromgxb_width NUMERIC "5"
-- Retrieval info: CONSTANT: reconfig_togxb_width NUMERIC "4"
-- Retrieval info: USED_PORT: busy 0 0 0 0 OUTPUT NODEFVAL "busy"
-- Retrieval info: USED_PORT: channel_reconfig_done 0 0 0 0 OUTPUT NODEFVAL "channel_reconfig_done"
-- Retrieval info: USED_PORT: error 0 0 0 0 OUTPUT NODEFVAL "error"
-- Retrieval info: USED_PORT: reconfig_address_en 0 0 0 0 OUTPUT NODEFVAL "reconfig_address_en"
-- Retrieval info: USED_PORT: reconfig_address_out 0 0 6 0 OUTPUT NODEFVAL "reconfig_address_out[5..0]"
-- Retrieval info: USED_PORT: reconfig_clk 0 0 0 0 INPUT NODEFVAL "reconfig_clk"
-- Retrieval info: USED_PORT: reconfig_data 0 0 16 0 INPUT NODEFVAL "reconfig_data[15..0]"
-- Retrieval info: USED_PORT: reconfig_fromgxb 0 0 5 0 INPUT NODEFVAL "reconfig_fromgxb[4..0]"
-- Retrieval info: USED_PORT: reconfig_reset 0 0 0 0 INPUT NODEFVAL "reconfig_reset"
-- Retrieval info: USED_PORT: reconfig_togxb 0 0 4 0 OUTPUT NODEFVAL "reconfig_togxb[3..0]"
-- Retrieval info: USED_PORT: write_all 0 0 0 0 INPUT NODEFVAL "write_all"
-- Retrieval info: CONNECT: @reconfig_clk 0 0 0 0 reconfig_clk 0 0 0 0
-- Retrieval info: CONNECT: @reconfig_data 0 0 16 0 reconfig_data 0 0 16 0
-- Retrieval info: CONNECT: @reconfig_fromgxb 0 0 5 0 reconfig_fromgxb 0 0 5 0
-- Retrieval info: CONNECT: @reconfig_mode_sel 0 0 1 1 GND 0 0 1 1
-- Retrieval info: CONNECT: @reconfig_mode_sel 0 0 1 2 GND 0 0 1 2
-- Retrieval info: CONNECT: @reconfig_mode_sel 0 0 1 0 VCC 0 0 1 0
-- Retrieval info: CONNECT: @reconfig_reset 0 0 0 0 reconfig_reset 0 0 0 0
-- Retrieval info: CONNECT: @write_all 0 0 0 0 write_all 0 0 0 0
-- Retrieval info: CONNECT: busy 0 0 0 0 @busy 0 0 0 0
-- Retrieval info: CONNECT: channel_reconfig_done 0 0 0 0 @channel_reconfig_done 0 0 0 0
-- Retrieval info: CONNECT: error 0 0 0 0 @error 0 0 0 0
-- Retrieval info: CONNECT: reconfig_address_en 0 0 0 0 @reconfig_address_en 0 0 0 0
-- Retrieval info: CONNECT: reconfig_address_out 0 0 6 0 @reconfig_address_out 0 0 6 0
-- Retrieval info: CONNECT: reconfig_togxb 0 0 4 0 @reconfig_togxb 0 0 4 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL ALTGX_RECONFIG_CIV.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL ALTGX_RECONFIG_CIV.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL ALTGX_RECONFIG_CIV.cmp TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL ALTGX_RECONFIG_CIV.bsf FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL ALTGX_RECONFIG_CIV_inst.vhd TRUE
-- Retrieval info: LIB_FILE: altera_mf
-- Retrieval info: LIB_FILE: lpm
